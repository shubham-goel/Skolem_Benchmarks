// Benchmark "ceiling32" written by ABC on Fri Sep 22 11:29:14 2017

module ceiling32 ( 
    \a[31] , \b[31] , \controllable_i[1] , \a[1] , \b[1] , \a[2] , \b[2] , \a[3] ,
    \b[3] , \a[4] , \b[4] , \a[5] , \b[5] , \a[6] , \b[6] , \a[7] , \b[7] ,
    \a[8] , \b[8] , \a[9] , \b[9] , \a[10] , \b[10] , \a[11] , \b[11] ,
    \a[12] , \b[12] , \a[13] , \b[13] , \a[14] , \b[14] , \a[15] , \b[15] ,
    \a[16] , \b[16] , \a[17] , \b[17] , \a[18] , \b[18] , \a[19] , \b[19] ,
    \a[20] , \b[20] , \a[21] , \b[21] , \a[22] , \b[22] , \a[23] , \b[23] ,
    \a[24] , \b[24] , \a[25] , \b[25] , \a[26] , \b[26] , \a[27] , \b[27] ,
    \a[28] , \b[28] , \a[29] , \b[29] , \a[30] , \b[30] , \a[0] , \b[0] ,
    \controllable_i[2] , \controllable_i[3] , \controllable_i[4] , \controllable_i[5] , \controllable_i[6] , \controllable_i[7] , \controllable_i[8] , \controllable_i[9] ,
    \controllable_i[10] , \controllable_i[11] , \controllable_i[12] , \controllable_i[13] , \controllable_i[14] , \controllable_i[15] , \controllable_i[16] , \controllable_i[17] ,
    \controllable_i[18] , \controllable_i[19] , \controllable_i[20] , \controllable_i[21] , \controllable_i[22] , \controllable_i[23] , \controllable_i[24] , \controllable_i[25] ,
    \controllable_i[26] , \controllable_i[27] , \controllable_i[28] , \controllable_i[29] , \controllable_i[30] , \controllable_i[31] ,
    n96  );
  input  \a[31] , \b[31] , \controllable_i[1] , \a[1] , \b[1] , \a[2] , \b[2] ,
    \a[3] , \b[3] , \a[4] , \b[4] , \a[5] , \b[5] , \a[6] , \b[6] , \a[7] ,
    \b[7] , \a[8] , \b[8] , \a[9] , \b[9] , \a[10] , \b[10] , \a[11] ,
    \b[11] , \a[12] , \b[12] , \a[13] , \b[13] , \a[14] , \b[14] , \a[15] ,
    \b[15] , \a[16] , \b[16] , \a[17] , \b[17] , \a[18] , \b[18] , \a[19] ,
    \b[19] , \a[20] , \b[20] , \a[21] , \b[21] , \a[22] , \b[22] , \a[23] ,
    \b[23] , \a[24] , \b[24] , \a[25] , \b[25] , \a[26] , \b[26] , \a[27] ,
    \b[27] , \a[28] , \b[28] , \a[29] , \b[29] , \a[30] , \b[30] , \a[0] ,
    \b[0] , \controllable_i[2] , \controllable_i[3] , \controllable_i[4] , \controllable_i[5] , \controllable_i[6] , \controllable_i[7] , \controllable_i[8] , \controllable_i[9] ,
    \controllable_i[10] , \controllable_i[11] , \controllable_i[12] , \controllable_i[13] , \controllable_i[14] , \controllable_i[15] , \controllable_i[16] , \controllable_i[17] ,
    \controllable_i[18] , \controllable_i[19] , \controllable_i[20] , \controllable_i[21] , \controllable_i[22] , \controllable_i[23] , \controllable_i[24] , \controllable_i[25] ,
    \controllable_i[26] , \controllable_i[27] , \controllable_i[28] , \controllable_i[29] , \controllable_i[30] , \controllable_i[31] ;
  output n96;
  wire n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656;
  assign n97 = \a[31]  & \b[31] ;
  assign n98 = ~\a[31]  & ~\b[31] ;
  assign n99 = ~n97 & ~n98;
  assign n100 = \a[1]  & \b[1] ;
  assign n101 = \a[2]  & \b[2] ;
  assign n102 = \a[3]  & \b[3] ;
  assign n103 = \a[4]  & \b[4] ;
  assign n104 = \a[5]  & \b[5] ;
  assign n105 = \a[6]  & \b[6] ;
  assign n106 = \a[7]  & \b[7] ;
  assign n107 = \a[8]  & \b[8] ;
  assign n108 = \a[9]  & \b[9] ;
  assign n109 = \a[10]  & \b[10] ;
  assign n110 = \a[11]  & \b[11] ;
  assign n111 = \a[12]  & \b[12] ;
  assign n112 = \a[13]  & \b[13] ;
  assign n113 = \a[14]  & \b[14] ;
  assign n114 = \a[15]  & \b[15] ;
  assign n115 = \a[16]  & \b[16] ;
  assign n116 = \a[17]  & \b[17] ;
  assign n117 = \a[18]  & \b[18] ;
  assign n118 = \a[19]  & \b[19] ;
  assign n119 = \a[20]  & \b[20] ;
  assign n120 = \a[21]  & \b[21] ;
  assign n121 = \a[22]  & \b[22] ;
  assign n122 = \a[23]  & \b[23] ;
  assign n123 = \a[24]  & \b[24] ;
  assign n124 = \a[25]  & \b[25] ;
  assign n125 = \a[26]  & \b[26] ;
  assign n126 = \a[27]  & \b[27] ;
  assign n127 = \a[28]  & \b[28] ;
  assign n128 = \a[29]  & \b[29] ;
  assign n129 = \a[30]  & \b[30] ;
  assign n130 = ~\a[30]  & ~\b[30] ;
  assign n131 = ~n129 & ~n130;
  assign n132 = n97 & n131;
  assign n133 = ~n129 & ~n132;
  assign n134 = ~\a[29]  & ~\b[29] ;
  assign n135 = ~n128 & ~n134;
  assign n136 = ~n133 & n135;
  assign n137 = ~n128 & ~n136;
  assign n138 = ~\a[28]  & ~\b[28] ;
  assign n139 = ~n127 & ~n138;
  assign n140 = ~n137 & n139;
  assign n141 = ~n127 & ~n140;
  assign n142 = ~\a[27]  & ~\b[27] ;
  assign n143 = ~n126 & ~n142;
  assign n144 = ~n141 & n143;
  assign n145 = ~n126 & ~n144;
  assign n146 = ~\a[26]  & ~\b[26] ;
  assign n147 = ~n125 & ~n146;
  assign n148 = ~n145 & n147;
  assign n149 = ~n125 & ~n148;
  assign n150 = ~\a[25]  & ~\b[25] ;
  assign n151 = ~n124 & ~n150;
  assign n152 = ~n149 & n151;
  assign n153 = ~n124 & ~n152;
  assign n154 = ~\a[24]  & ~\b[24] ;
  assign n155 = ~n123 & ~n154;
  assign n156 = ~n153 & n155;
  assign n157 = ~n123 & ~n156;
  assign n158 = ~\a[23]  & ~\b[23] ;
  assign n159 = ~n122 & ~n158;
  assign n160 = ~n157 & n159;
  assign n161 = ~n122 & ~n160;
  assign n162 = ~\a[22]  & ~\b[22] ;
  assign n163 = ~n121 & ~n162;
  assign n164 = ~n161 & n163;
  assign n165 = ~n121 & ~n164;
  assign n166 = ~\a[21]  & ~\b[21] ;
  assign n167 = ~n120 & ~n166;
  assign n168 = ~n165 & n167;
  assign n169 = ~n120 & ~n168;
  assign n170 = ~\a[20]  & ~\b[20] ;
  assign n171 = ~n119 & ~n170;
  assign n172 = ~n169 & n171;
  assign n173 = ~n119 & ~n172;
  assign n174 = ~\a[19]  & ~\b[19] ;
  assign n175 = ~n118 & ~n174;
  assign n176 = ~n173 & n175;
  assign n177 = ~n118 & ~n176;
  assign n178 = ~\a[18]  & ~\b[18] ;
  assign n179 = ~n117 & ~n178;
  assign n180 = ~n177 & n179;
  assign n181 = ~n117 & ~n180;
  assign n182 = ~\a[17]  & ~\b[17] ;
  assign n183 = ~n116 & ~n182;
  assign n184 = ~n181 & n183;
  assign n185 = ~n116 & ~n184;
  assign n186 = ~\a[16]  & ~\b[16] ;
  assign n187 = ~n115 & ~n186;
  assign n188 = ~n185 & n187;
  assign n189 = ~n115 & ~n188;
  assign n190 = ~\a[15]  & ~\b[15] ;
  assign n191 = ~n114 & ~n190;
  assign n192 = ~n189 & n191;
  assign n193 = ~n114 & ~n192;
  assign n194 = ~\a[14]  & ~\b[14] ;
  assign n195 = ~n113 & ~n194;
  assign n196 = ~n193 & n195;
  assign n197 = ~n113 & ~n196;
  assign n198 = ~\a[13]  & ~\b[13] ;
  assign n199 = ~n112 & ~n198;
  assign n200 = ~n197 & n199;
  assign n201 = ~n112 & ~n200;
  assign n202 = ~\a[12]  & ~\b[12] ;
  assign n203 = ~n111 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = ~n111 & ~n204;
  assign n206 = ~\a[11]  & ~\b[11] ;
  assign n207 = ~n110 & ~n206;
  assign n208 = ~n205 & n207;
  assign n209 = ~n110 & ~n208;
  assign n210 = ~\a[10]  & ~\b[10] ;
  assign n211 = ~n109 & ~n210;
  assign n212 = ~n209 & n211;
  assign n213 = ~n109 & ~n212;
  assign n214 = ~\a[9]  & ~\b[9] ;
  assign n215 = ~n108 & ~n214;
  assign n216 = ~n213 & n215;
  assign n217 = ~n108 & ~n216;
  assign n218 = ~\a[8]  & ~\b[8] ;
  assign n219 = ~n107 & ~n218;
  assign n220 = ~n217 & n219;
  assign n221 = ~n107 & ~n220;
  assign n222 = ~\a[7]  & ~\b[7] ;
  assign n223 = ~n106 & ~n222;
  assign n224 = ~n221 & n223;
  assign n225 = ~n106 & ~n224;
  assign n226 = ~\a[6]  & ~\b[6] ;
  assign n227 = ~n105 & ~n226;
  assign n228 = ~n225 & n227;
  assign n229 = ~n105 & ~n228;
  assign n230 = ~\a[5]  & ~\b[5] ;
  assign n231 = ~n104 & ~n230;
  assign n232 = ~n229 & n231;
  assign n233 = ~n104 & ~n232;
  assign n234 = ~\a[4]  & ~\b[4] ;
  assign n235 = ~n103 & ~n234;
  assign n236 = ~n233 & n235;
  assign n237 = ~n103 & ~n236;
  assign n238 = ~\a[3]  & ~\b[3] ;
  assign n239 = ~n102 & ~n238;
  assign n240 = ~n237 & n239;
  assign n241 = ~n102 & ~n240;
  assign n242 = ~\a[2]  & ~\b[2] ;
  assign n243 = ~n101 & ~n242;
  assign n244 = ~n241 & n243;
  assign n245 = ~n101 & ~n244;
  assign n246 = ~\a[1]  & ~\b[1] ;
  assign n247 = ~n100 & ~n246;
  assign n248 = ~n245 & n247;
  assign n249 = ~n100 & ~n248;
  assign n250 = \a[0]  & \b[0] ;
  assign n251 = ~\a[0]  & ~\b[0] ;
  assign n252 = ~n250 & ~n251;
  assign n253 = ~n249 & n252;
  assign n254 = n249 & ~n252;
  assign n255 = ~n253 & ~n254;
  assign n256 = \controllable_i[1]  & ~n255;
  assign n257 = ~\controllable_i[1]  & n255;
  assign n258 = ~n256 & ~n257;
  assign n259 = n245 & ~n247;
  assign n260 = ~n248 & ~n259;
  assign n261 = \controllable_i[2]  & ~n260;
  assign n262 = ~\controllable_i[2]  & n260;
  assign n263 = ~n261 & ~n262;
  assign n264 = n258 & n263;
  assign n265 = n241 & ~n243;
  assign n266 = ~n244 & ~n265;
  assign n267 = \controllable_i[3]  & ~n266;
  assign n268 = ~\controllable_i[3]  & n266;
  assign n269 = ~n267 & ~n268;
  assign n270 = n264 & n269;
  assign n271 = n237 & ~n239;
  assign n272 = ~n240 & ~n271;
  assign n273 = \controllable_i[4]  & ~n272;
  assign n274 = ~\controllable_i[4]  & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = n270 & n275;
  assign n277 = n233 & ~n235;
  assign n278 = ~n236 & ~n277;
  assign n279 = \controllable_i[5]  & ~n278;
  assign n280 = ~\controllable_i[5]  & n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = n276 & n281;
  assign n283 = n229 & ~n231;
  assign n284 = ~n232 & ~n283;
  assign n285 = \controllable_i[6]  & ~n284;
  assign n286 = ~\controllable_i[6]  & n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = n282 & n287;
  assign n289 = n225 & ~n227;
  assign n290 = ~n228 & ~n289;
  assign n291 = \controllable_i[7]  & ~n290;
  assign n292 = ~\controllable_i[7]  & n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = n288 & n293;
  assign n295 = n221 & ~n223;
  assign n296 = ~n224 & ~n295;
  assign n297 = \controllable_i[8]  & ~n296;
  assign n298 = ~\controllable_i[8]  & n296;
  assign n299 = ~n297 & ~n298;
  assign n300 = n294 & n299;
  assign n301 = n217 & ~n219;
  assign n302 = ~n220 & ~n301;
  assign n303 = \controllable_i[9]  & ~n302;
  assign n304 = ~\controllable_i[9]  & n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = n300 & n305;
  assign n307 = n213 & ~n215;
  assign n308 = ~n216 & ~n307;
  assign n309 = \controllable_i[10]  & ~n308;
  assign n310 = ~\controllable_i[10]  & n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = n306 & n311;
  assign n313 = n209 & ~n211;
  assign n314 = ~n212 & ~n313;
  assign n315 = \controllable_i[11]  & ~n314;
  assign n316 = ~\controllable_i[11]  & n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = n312 & n317;
  assign n319 = n205 & ~n207;
  assign n320 = ~n208 & ~n319;
  assign n321 = \controllable_i[12]  & ~n320;
  assign n322 = ~\controllable_i[12]  & n320;
  assign n323 = ~n321 & ~n322;
  assign n324 = n318 & n323;
  assign n325 = n201 & ~n203;
  assign n326 = ~n204 & ~n325;
  assign n327 = \controllable_i[13]  & ~n326;
  assign n328 = ~\controllable_i[13]  & n326;
  assign n329 = ~n327 & ~n328;
  assign n330 = n324 & n329;
  assign n331 = n197 & ~n199;
  assign n332 = ~n200 & ~n331;
  assign n333 = \controllable_i[14]  & ~n332;
  assign n334 = ~\controllable_i[14]  & n332;
  assign n335 = ~n333 & ~n334;
  assign n336 = n330 & n335;
  assign n337 = n193 & ~n195;
  assign n338 = ~n196 & ~n337;
  assign n339 = \controllable_i[15]  & ~n338;
  assign n340 = ~\controllable_i[15]  & n338;
  assign n341 = ~n339 & ~n340;
  assign n342 = n336 & n341;
  assign n343 = n189 & ~n191;
  assign n344 = ~n192 & ~n343;
  assign n345 = \controllable_i[16]  & ~n344;
  assign n346 = ~\controllable_i[16]  & n344;
  assign n347 = ~n345 & ~n346;
  assign n348 = n342 & n347;
  assign n349 = n185 & ~n187;
  assign n350 = ~n188 & ~n349;
  assign n351 = \controllable_i[17]  & ~n350;
  assign n352 = ~\controllable_i[17]  & n350;
  assign n353 = ~n351 & ~n352;
  assign n354 = n348 & n353;
  assign n355 = n181 & ~n183;
  assign n356 = ~n184 & ~n355;
  assign n357 = \controllable_i[18]  & ~n356;
  assign n358 = ~\controllable_i[18]  & n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = n354 & n359;
  assign n361 = n177 & ~n179;
  assign n362 = ~n180 & ~n361;
  assign n363 = \controllable_i[19]  & ~n362;
  assign n364 = ~\controllable_i[19]  & n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = n360 & n365;
  assign n367 = n173 & ~n175;
  assign n368 = ~n176 & ~n367;
  assign n369 = \controllable_i[20]  & ~n368;
  assign n370 = ~\controllable_i[20]  & n368;
  assign n371 = ~n369 & ~n370;
  assign n372 = n366 & n371;
  assign n373 = n169 & ~n171;
  assign n374 = ~n172 & ~n373;
  assign n375 = \controllable_i[21]  & ~n374;
  assign n376 = ~\controllable_i[21]  & n374;
  assign n377 = ~n375 & ~n376;
  assign n378 = n372 & n377;
  assign n379 = n165 & ~n167;
  assign n380 = ~n168 & ~n379;
  assign n381 = \controllable_i[22]  & ~n380;
  assign n382 = ~\controllable_i[22]  & n380;
  assign n383 = ~n381 & ~n382;
  assign n384 = n378 & n383;
  assign n385 = n161 & ~n163;
  assign n386 = ~n164 & ~n385;
  assign n387 = \controllable_i[23]  & ~n386;
  assign n388 = ~\controllable_i[23]  & n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = n384 & n389;
  assign n391 = n157 & ~n159;
  assign n392 = ~n160 & ~n391;
  assign n393 = \controllable_i[24]  & ~n392;
  assign n394 = ~\controllable_i[24]  & n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = n390 & n395;
  assign n397 = n153 & ~n155;
  assign n398 = ~n156 & ~n397;
  assign n399 = \controllable_i[25]  & ~n398;
  assign n400 = ~\controllable_i[25]  & n398;
  assign n401 = ~n399 & ~n400;
  assign n402 = n396 & n401;
  assign n403 = n149 & ~n151;
  assign n404 = ~n152 & ~n403;
  assign n405 = \controllable_i[26]  & ~n404;
  assign n406 = ~\controllable_i[26]  & n404;
  assign n407 = ~n405 & ~n406;
  assign n408 = n402 & n407;
  assign n409 = n145 & ~n147;
  assign n410 = ~n148 & ~n409;
  assign n411 = \controllable_i[27]  & ~n410;
  assign n412 = ~\controllable_i[27]  & n410;
  assign n413 = ~n411 & ~n412;
  assign n414 = n408 & n413;
  assign n415 = n141 & ~n143;
  assign n416 = ~n144 & ~n415;
  assign n417 = \controllable_i[28]  & ~n416;
  assign n418 = ~\controllable_i[28]  & n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = n414 & n419;
  assign n421 = n137 & ~n139;
  assign n422 = ~n140 & ~n421;
  assign n423 = \controllable_i[29]  & ~n422;
  assign n424 = ~\controllable_i[29]  & n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = n420 & n425;
  assign n427 = n133 & ~n135;
  assign n428 = ~n136 & ~n427;
  assign n429 = \controllable_i[30]  & ~n428;
  assign n430 = ~\controllable_i[30]  & n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = n426 & n431;
  assign n433 = ~n97 & ~n131;
  assign n434 = ~n132 & ~n433;
  assign n435 = \controllable_i[31]  & ~n434;
  assign n436 = ~\controllable_i[31]  & n434;
  assign n437 = ~n435 & ~n436;
  assign n438 = n432 & n437;
  assign n439 = ~n99 & n438;
  assign n440 = n99 & n434;
  assign n441 = n428 & n440;
  assign n442 = n422 & n441;
  assign n443 = n416 & n442;
  assign n444 = n410 & n443;
  assign n445 = n404 & n444;
  assign n446 = n398 & n445;
  assign n447 = n392 & n446;
  assign n448 = n386 & n447;
  assign n449 = n380 & n448;
  assign n450 = n374 & n449;
  assign n451 = n368 & n450;
  assign n452 = n362 & n451;
  assign n453 = n356 & n452;
  assign n454 = n350 & n453;
  assign n455 = n344 & n454;
  assign n456 = n338 & n455;
  assign n457 = n332 & n456;
  assign n458 = n326 & n457;
  assign n459 = n320 & n458;
  assign n460 = n314 & n459;
  assign n461 = n308 & n460;
  assign n462 = n302 & n461;
  assign n463 = n296 & n462;
  assign n464 = n290 & n463;
  assign n465 = n284 & n464;
  assign n466 = n278 & n465;
  assign n467 = n272 & n466;
  assign n468 = n266 & n467;
  assign n469 = n260 & n468;
  assign n470 = n255 & n469;
  assign n471 = ~n255 & ~n469;
  assign n472 = ~n470 & ~n471;
  assign n473 = \controllable_i[1]  & ~n472;
  assign n474 = ~\controllable_i[1]  & n472;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n260 & ~n468;
  assign n477 = ~n469 & ~n476;
  assign n478 = \controllable_i[2]  & ~n477;
  assign n479 = ~\controllable_i[2]  & n477;
  assign n480 = ~n478 & ~n479;
  assign n481 = n475 & n480;
  assign n482 = ~n266 & ~n467;
  assign n483 = ~n468 & ~n482;
  assign n484 = \controllable_i[3]  & ~n483;
  assign n485 = ~\controllable_i[3]  & n483;
  assign n486 = ~n484 & ~n485;
  assign n487 = n481 & n486;
  assign n488 = ~n272 & ~n466;
  assign n489 = ~n467 & ~n488;
  assign n490 = \controllable_i[4]  & ~n489;
  assign n491 = ~\controllable_i[4]  & n489;
  assign n492 = ~n490 & ~n491;
  assign n493 = n487 & n492;
  assign n494 = ~n278 & ~n465;
  assign n495 = ~n466 & ~n494;
  assign n496 = \controllable_i[5]  & ~n495;
  assign n497 = ~\controllable_i[5]  & n495;
  assign n498 = ~n496 & ~n497;
  assign n499 = n493 & n498;
  assign n500 = ~n284 & ~n464;
  assign n501 = ~n465 & ~n500;
  assign n502 = \controllable_i[6]  & ~n501;
  assign n503 = ~\controllable_i[6]  & n501;
  assign n504 = ~n502 & ~n503;
  assign n505 = n499 & n504;
  assign n506 = ~n290 & ~n463;
  assign n507 = ~n464 & ~n506;
  assign n508 = \controllable_i[7]  & ~n507;
  assign n509 = ~\controllable_i[7]  & n507;
  assign n510 = ~n508 & ~n509;
  assign n511 = n505 & n510;
  assign n512 = ~n296 & ~n462;
  assign n513 = ~n463 & ~n512;
  assign n514 = \controllable_i[8]  & ~n513;
  assign n515 = ~\controllable_i[8]  & n513;
  assign n516 = ~n514 & ~n515;
  assign n517 = n511 & n516;
  assign n518 = ~n302 & ~n461;
  assign n519 = ~n462 & ~n518;
  assign n520 = \controllable_i[9]  & ~n519;
  assign n521 = ~\controllable_i[9]  & n519;
  assign n522 = ~n520 & ~n521;
  assign n523 = n517 & n522;
  assign n524 = ~n308 & ~n460;
  assign n525 = ~n461 & ~n524;
  assign n526 = \controllable_i[10]  & ~n525;
  assign n527 = ~\controllable_i[10]  & n525;
  assign n528 = ~n526 & ~n527;
  assign n529 = n523 & n528;
  assign n530 = ~n314 & ~n459;
  assign n531 = ~n460 & ~n530;
  assign n532 = \controllable_i[11]  & ~n531;
  assign n533 = ~\controllable_i[11]  & n531;
  assign n534 = ~n532 & ~n533;
  assign n535 = n529 & n534;
  assign n536 = ~n320 & ~n458;
  assign n537 = ~n459 & ~n536;
  assign n538 = \controllable_i[12]  & ~n537;
  assign n539 = ~\controllable_i[12]  & n537;
  assign n540 = ~n538 & ~n539;
  assign n541 = n535 & n540;
  assign n542 = ~n326 & ~n457;
  assign n543 = ~n458 & ~n542;
  assign n544 = \controllable_i[13]  & ~n543;
  assign n545 = ~\controllable_i[13]  & n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = n541 & n546;
  assign n548 = ~n332 & ~n456;
  assign n549 = ~n457 & ~n548;
  assign n550 = \controllable_i[14]  & ~n549;
  assign n551 = ~\controllable_i[14]  & n549;
  assign n552 = ~n550 & ~n551;
  assign n553 = n547 & n552;
  assign n554 = ~n338 & ~n455;
  assign n555 = ~n456 & ~n554;
  assign n556 = \controllable_i[15]  & ~n555;
  assign n557 = ~\controllable_i[15]  & n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = n553 & n558;
  assign n560 = ~n344 & ~n454;
  assign n561 = ~n455 & ~n560;
  assign n562 = \controllable_i[16]  & ~n561;
  assign n563 = ~\controllable_i[16]  & n561;
  assign n564 = ~n562 & ~n563;
  assign n565 = n559 & n564;
  assign n566 = ~n350 & ~n453;
  assign n567 = ~n454 & ~n566;
  assign n568 = \controllable_i[17]  & ~n567;
  assign n569 = ~\controllable_i[17]  & n567;
  assign n570 = ~n568 & ~n569;
  assign n571 = n565 & n570;
  assign n572 = ~n356 & ~n452;
  assign n573 = ~n453 & ~n572;
  assign n574 = \controllable_i[18]  & ~n573;
  assign n575 = ~\controllable_i[18]  & n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = n571 & n576;
  assign n578 = ~n362 & ~n451;
  assign n579 = ~n452 & ~n578;
  assign n580 = \controllable_i[19]  & ~n579;
  assign n581 = ~\controllable_i[19]  & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = n577 & n582;
  assign n584 = ~n368 & ~n450;
  assign n585 = ~n451 & ~n584;
  assign n586 = \controllable_i[20]  & ~n585;
  assign n587 = ~\controllable_i[20]  & n585;
  assign n588 = ~n586 & ~n587;
  assign n589 = n583 & n588;
  assign n590 = ~n374 & ~n449;
  assign n591 = ~n450 & ~n590;
  assign n592 = \controllable_i[21]  & ~n591;
  assign n593 = ~\controllable_i[21]  & n591;
  assign n594 = ~n592 & ~n593;
  assign n595 = n589 & n594;
  assign n596 = ~n380 & ~n448;
  assign n597 = ~n449 & ~n596;
  assign n598 = \controllable_i[22]  & ~n597;
  assign n599 = ~\controllable_i[22]  & n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = n595 & n600;
  assign n602 = ~n386 & ~n447;
  assign n603 = ~n448 & ~n602;
  assign n604 = \controllable_i[23]  & ~n603;
  assign n605 = ~\controllable_i[23]  & n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = n601 & n606;
  assign n608 = ~n392 & ~n446;
  assign n609 = ~n447 & ~n608;
  assign n610 = \controllable_i[24]  & ~n609;
  assign n611 = ~\controllable_i[24]  & n609;
  assign n612 = ~n610 & ~n611;
  assign n613 = n607 & n612;
  assign n614 = ~n398 & ~n445;
  assign n615 = ~n446 & ~n614;
  assign n616 = \controllable_i[25]  & ~n615;
  assign n617 = ~\controllable_i[25]  & n615;
  assign n618 = ~n616 & ~n617;
  assign n619 = n613 & n618;
  assign n620 = ~n404 & ~n444;
  assign n621 = ~n445 & ~n620;
  assign n622 = \controllable_i[26]  & ~n621;
  assign n623 = ~\controllable_i[26]  & n621;
  assign n624 = ~n622 & ~n623;
  assign n625 = n619 & n624;
  assign n626 = ~n410 & ~n443;
  assign n627 = ~n444 & ~n626;
  assign n628 = \controllable_i[27]  & ~n627;
  assign n629 = ~\controllable_i[27]  & n627;
  assign n630 = ~n628 & ~n629;
  assign n631 = n625 & n630;
  assign n632 = ~n416 & ~n442;
  assign n633 = ~n443 & ~n632;
  assign n634 = \controllable_i[28]  & ~n633;
  assign n635 = ~\controllable_i[28]  & n633;
  assign n636 = ~n634 & ~n635;
  assign n637 = n631 & n636;
  assign n638 = ~n422 & ~n441;
  assign n639 = ~n442 & ~n638;
  assign n640 = \controllable_i[29]  & ~n639;
  assign n641 = ~\controllable_i[29]  & n639;
  assign n642 = ~n640 & ~n641;
  assign n643 = n637 & n642;
  assign n644 = ~n428 & ~n440;
  assign n645 = ~n441 & ~n644;
  assign n646 = \controllable_i[30]  & ~n645;
  assign n647 = ~\controllable_i[30]  & n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = n643 & n648;
  assign n650 = ~n99 & ~n434;
  assign n651 = ~n440 & ~n650;
  assign n652 = \controllable_i[31]  & ~n651;
  assign n653 = ~\controllable_i[31]  & n651;
  assign n654 = ~n652 & ~n653;
  assign n655 = n649 & n654;
  assign n656 = n99 & n655;
  assign n96 = n439 | n656;
endmodule


