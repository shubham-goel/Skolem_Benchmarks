// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module factorization20_simplified ( i2[19], i2[18], i2[17], i2[16], i2[15], i2[14], i2[13], i2[12], i2[11], i2[10], i1[19], i1[18], i1[17], i1[16], i1[15], i1[14], i1[13], i1[12], i1[11], i1[10], a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], o_1 );
input i2[19];
input i2[18];
input i2[17];
input i2[16];
input i2[15];
input i2[14];
input i2[13];
input i2[12];
input i2[11];
input i2[10];
input i1[19];
input i1[18];
input i1[17];
input i1[16];
input i1[15];
input i1[14];
input i1[13];
input i1[12];
input i1[11];
input i1[10];
input a[0];
input a[1];
input a[2];
input a[3];
input a[4];
input a[5];
input a[6];
input a[7];
input a[8];
input a[9];
input a[10];
input a[11];
input a[12];
input a[13];
input a[14];
input a[15];
input a[16];
input a[17];
input a[18];
input a[19];
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
assign n_1 =  i2[10] &  i1[10];
assign n_2 =  i2[10] &  i1[11];
assign n_3 =  i2[10] &  i1[12];
assign n_4 =  i2[10] &  i1[13];
assign n_5 =  i2[10] &  i1[14];
assign n_6 =  i2[10] &  i1[15];
assign n_7 =  i2[10] &  i1[16];
assign n_8 =  i2[10] &  i1[17];
assign n_9 =  i2[11] &  i1[18];
assign n_10 =  i2[10] &  i1[19];
assign n_11 =  n_9 &  n_10;
assign n_12 =  i2[12] &  i1[18];
assign n_13 =  i2[11] &  i1[19];
assign n_14 =  n_12 &  n_13;
assign n_15 =  i2[13] &  i1[18];
assign n_16 =  i2[12] &  i1[19];
assign n_17 =  n_15 &  n_16;
assign n_18 =  i2[14] &  i1[18];
assign n_19 =  i2[13] &  i1[19];
assign n_20 =  n_18 &  n_19;
assign n_21 =  i2[15] &  i1[18];
assign n_22 =  i2[14] &  i1[19];
assign n_23 =  n_21 &  n_22;
assign n_24 =  i2[16] &  i1[18];
assign n_25 =  i2[15] &  i1[19];
assign n_26 =  n_24 &  n_25;
assign n_27 =  i2[17] &  i1[18];
assign n_28 =  i2[16] &  i1[19];
assign n_29 =  n_27 &  n_28;
assign n_30 =  i2[18] &  i1[19];
assign n_31 =  i2[19] &  i1[18];
assign n_32 =  n_30 &  n_31;
assign n_33 =  i2[18] &  i1[18];
assign n_34 =  i2[17] &  i1[19];
assign n_35 =  n_33 &  n_34;
assign n_36 = ~n_32 & ~n_35;
assign n_37 = ~n_27 & ~n_28;
assign n_38 = ~n_37 & ~n_29;
assign n_39 = ~n_36 &  n_38;
assign n_40 = ~n_29 & ~n_39;
assign n_41 = ~n_24 & ~n_25;
assign n_42 = ~n_41 & ~n_26;
assign n_43 = ~n_40 &  n_42;
assign n_44 = ~n_26 & ~n_43;
assign n_45 = ~n_21 & ~n_22;
assign n_46 = ~n_45 & ~n_23;
assign n_47 = ~n_44 &  n_46;
assign n_48 = ~n_23 & ~n_47;
assign n_49 = ~n_18 & ~n_19;
assign n_50 = ~n_49 & ~n_20;
assign n_51 = ~n_48 &  n_50;
assign n_52 = ~n_20 & ~n_51;
assign n_53 = ~n_15 & ~n_16;
assign n_54 = ~n_53 & ~n_17;
assign n_55 = ~n_52 &  n_54;
assign n_56 = ~n_17 & ~n_55;
assign n_57 = ~n_12 & ~n_13;
assign n_58 = ~n_57 & ~n_14;
assign n_59 = ~n_56 &  n_58;
assign n_60 = ~n_14 & ~n_59;
assign n_61 = ~n_9 & ~n_10;
assign n_62 = ~n_61 & ~n_11;
assign n_63 = ~n_60 &  n_62;
assign n_64 = ~n_11 & ~n_63;
assign n_65 =  i2[10] &  i1[18];
assign n_66 = ~n_64 &  n_65;
assign n_67 =  n_8 &  n_66;
assign n_68 =  i2[11] &  i1[17];
assign n_69 =  n_64 & ~n_65;
assign n_70 = ~n_66 & ~n_69;
assign n_71 =  n_68 &  n_70;
assign n_72 =  n_60 & ~n_62;
assign n_73 = ~n_63 & ~n_72;
assign n_74 =  i2[12] &  i1[17];
assign n_75 =  n_73 &  n_74;
assign n_76 =  n_56 & ~n_58;
assign n_77 = ~n_59 & ~n_76;
assign n_78 =  i2[13] &  i1[17];
assign n_79 =  n_77 &  n_78;
assign n_80 =  n_52 & ~n_54;
assign n_81 = ~n_55 & ~n_80;
assign n_82 =  i2[14] &  i1[17];
assign n_83 =  n_81 &  n_82;
assign n_84 =  n_48 & ~n_50;
assign n_85 = ~n_51 & ~n_84;
assign n_86 =  i2[15] &  i1[17];
assign n_87 =  n_85 &  n_86;
assign n_88 =  n_44 & ~n_46;
assign n_89 = ~n_47 & ~n_88;
assign n_90 =  i2[16] &  i1[17];
assign n_91 =  n_89 &  n_90;
assign n_92 =  n_40 & ~n_42;
assign n_93 = ~n_43 & ~n_92;
assign n_94 =  i2[17] &  i1[17];
assign n_95 =  n_93 &  n_94;
assign n_96 =  n_36 & ~n_38;
assign n_97 = ~n_39 & ~n_96;
assign n_98 =  i2[18] &  i1[17];
assign n_99 =  n_97 &  n_98;
assign n_100 =  i2[19] &  i1[17];
assign n_101 =  n_32 &  n_35;
assign n_102 = ~n_36 & ~n_101;
assign n_103 = ~n_33 & ~n_34;
assign n_104 = ~n_102 & ~n_103;
assign n_105 =  n_100 &  n_104;
assign n_106 = ~n_97 & ~n_98;
assign n_107 = ~n_99 & ~n_106;
assign n_108 =  n_105 &  n_107;
assign n_109 = ~n_99 & ~n_108;
assign n_110 = ~n_93 & ~n_94;
assign n_111 = ~n_95 & ~n_110;
assign n_112 = ~n_109 &  n_111;
assign n_113 = ~n_95 & ~n_112;
assign n_114 = ~n_89 & ~n_90;
assign n_115 = ~n_91 & ~n_114;
assign n_116 = ~n_113 &  n_115;
assign n_117 = ~n_91 & ~n_116;
assign n_118 = ~n_85 & ~n_86;
assign n_119 = ~n_87 & ~n_118;
assign n_120 = ~n_117 &  n_119;
assign n_121 = ~n_87 & ~n_120;
assign n_122 = ~n_81 & ~n_82;
assign n_123 = ~n_83 & ~n_122;
assign n_124 = ~n_121 &  n_123;
assign n_125 = ~n_83 & ~n_124;
assign n_126 = ~n_77 & ~n_78;
assign n_127 = ~n_79 & ~n_126;
assign n_128 = ~n_125 &  n_127;
assign n_129 = ~n_79 & ~n_128;
assign n_130 = ~n_73 & ~n_74;
assign n_131 = ~n_75 & ~n_130;
assign n_132 = ~n_129 &  n_131;
assign n_133 = ~n_75 & ~n_132;
assign n_134 = ~n_68 & ~n_70;
assign n_135 = ~n_71 & ~n_134;
assign n_136 = ~n_133 &  n_135;
assign n_137 = ~n_71 & ~n_136;
assign n_138 = ~n_8 & ~n_66;
assign n_139 = ~n_67 & ~n_138;
assign n_140 = ~n_137 &  n_139;
assign n_141 = ~n_67 & ~n_140;
assign n_142 =  n_7 & ~n_141;
assign n_143 =  i2[11] &  i1[16];
assign n_144 =  n_137 & ~n_139;
assign n_145 = ~n_140 & ~n_144;
assign n_146 =  n_143 &  n_145;
assign n_147 =  i2[12] &  i1[16];
assign n_148 =  n_133 & ~n_135;
assign n_149 = ~n_136 & ~n_148;
assign n_150 =  n_147 &  n_149;
assign n_151 =  n_129 & ~n_131;
assign n_152 = ~n_132 & ~n_151;
assign n_153 =  i2[13] &  i1[16];
assign n_154 =  n_152 &  n_153;
assign n_155 =  n_125 & ~n_127;
assign n_156 = ~n_128 & ~n_155;
assign n_157 =  i2[14] &  i1[16];
assign n_158 =  n_156 &  n_157;
assign n_159 =  n_121 & ~n_123;
assign n_160 = ~n_124 & ~n_159;
assign n_161 =  i2[15] &  i1[16];
assign n_162 =  n_160 &  n_161;
assign n_163 =  n_117 & ~n_119;
assign n_164 = ~n_120 & ~n_163;
assign n_165 =  i2[16] &  i1[16];
assign n_166 =  n_164 &  n_165;
assign n_167 =  n_113 & ~n_115;
assign n_168 = ~n_116 & ~n_167;
assign n_169 =  i2[17] &  i1[16];
assign n_170 =  n_168 &  n_169;
assign n_171 =  n_109 & ~n_111;
assign n_172 = ~n_112 & ~n_171;
assign n_173 =  i2[18] &  i1[16];
assign n_174 =  n_172 &  n_173;
assign n_175 = ~n_105 & ~n_107;
assign n_176 = ~n_108 & ~n_175;
assign n_177 =  i2[19] &  i1[16];
assign n_178 =  n_176 &  n_177;
assign n_179 = ~n_172 & ~n_173;
assign n_180 = ~n_174 & ~n_179;
assign n_181 =  n_178 &  n_180;
assign n_182 = ~n_174 & ~n_181;
assign n_183 = ~n_168 & ~n_169;
assign n_184 = ~n_170 & ~n_183;
assign n_185 = ~n_182 &  n_184;
assign n_186 = ~n_170 & ~n_185;
assign n_187 = ~n_164 & ~n_165;
assign n_188 = ~n_166 & ~n_187;
assign n_189 = ~n_186 &  n_188;
assign n_190 = ~n_166 & ~n_189;
assign n_191 = ~n_160 & ~n_161;
assign n_192 = ~n_162 & ~n_191;
assign n_193 = ~n_190 &  n_192;
assign n_194 = ~n_162 & ~n_193;
assign n_195 = ~n_156 & ~n_157;
assign n_196 = ~n_158 & ~n_195;
assign n_197 = ~n_194 &  n_196;
assign n_198 = ~n_158 & ~n_197;
assign n_199 = ~n_152 & ~n_153;
assign n_200 = ~n_154 & ~n_199;
assign n_201 = ~n_198 &  n_200;
assign n_202 = ~n_154 & ~n_201;
assign n_203 = ~n_147 & ~n_149;
assign n_204 = ~n_150 & ~n_203;
assign n_205 = ~n_202 &  n_204;
assign n_206 = ~n_150 & ~n_205;
assign n_207 = ~n_143 & ~n_145;
assign n_208 = ~n_146 & ~n_207;
assign n_209 = ~n_206 &  n_208;
assign n_210 = ~n_146 & ~n_209;
assign n_211 = ~n_7 &  n_141;
assign n_212 = ~n_142 & ~n_211;
assign n_213 = ~n_210 &  n_212;
assign n_214 = ~n_142 & ~n_213;
assign n_215 =  n_6 & ~n_214;
assign n_216 =  i2[11] &  i1[15];
assign n_217 =  n_210 & ~n_212;
assign n_218 = ~n_213 & ~n_217;
assign n_219 =  n_216 &  n_218;
assign n_220 =  i2[12] &  i1[15];
assign n_221 =  n_206 & ~n_208;
assign n_222 = ~n_209 & ~n_221;
assign n_223 =  n_220 &  n_222;
assign n_224 =  i2[13] &  i1[15];
assign n_225 =  n_202 & ~n_204;
assign n_226 = ~n_205 & ~n_225;
assign n_227 =  n_224 &  n_226;
assign n_228 =  n_198 & ~n_200;
assign n_229 = ~n_201 & ~n_228;
assign n_230 =  i2[14] &  i1[15];
assign n_231 =  n_229 &  n_230;
assign n_232 =  n_194 & ~n_196;
assign n_233 = ~n_197 & ~n_232;
assign n_234 =  i2[15] &  i1[15];
assign n_235 =  n_233 &  n_234;
assign n_236 =  n_190 & ~n_192;
assign n_237 = ~n_193 & ~n_236;
assign n_238 =  i2[16] &  i1[15];
assign n_239 =  n_237 &  n_238;
assign n_240 =  n_186 & ~n_188;
assign n_241 = ~n_189 & ~n_240;
assign n_242 =  i2[17] &  i1[15];
assign n_243 =  n_241 &  n_242;
assign n_244 =  n_182 & ~n_184;
assign n_245 = ~n_185 & ~n_244;
assign n_246 =  i2[18] &  i1[15];
assign n_247 =  n_245 &  n_246;
assign n_248 = ~n_178 & ~n_180;
assign n_249 = ~n_181 & ~n_248;
assign n_250 =  i2[19] &  i1[15];
assign n_251 =  n_249 &  n_250;
assign n_252 = ~n_245 & ~n_246;
assign n_253 = ~n_247 & ~n_252;
assign n_254 =  n_251 &  n_253;
assign n_255 = ~n_247 & ~n_254;
assign n_256 = ~n_241 & ~n_242;
assign n_257 = ~n_243 & ~n_256;
assign n_258 = ~n_255 &  n_257;
assign n_259 = ~n_243 & ~n_258;
assign n_260 = ~n_237 & ~n_238;
assign n_261 = ~n_239 & ~n_260;
assign n_262 = ~n_259 &  n_261;
assign n_263 = ~n_239 & ~n_262;
assign n_264 = ~n_233 & ~n_234;
assign n_265 = ~n_235 & ~n_264;
assign n_266 = ~n_263 &  n_265;
assign n_267 = ~n_235 & ~n_266;
assign n_268 = ~n_229 & ~n_230;
assign n_269 = ~n_231 & ~n_268;
assign n_270 = ~n_267 &  n_269;
assign n_271 = ~n_231 & ~n_270;
assign n_272 = ~n_224 & ~n_226;
assign n_273 = ~n_227 & ~n_272;
assign n_274 = ~n_271 &  n_273;
assign n_275 = ~n_227 & ~n_274;
assign n_276 = ~n_220 & ~n_222;
assign n_277 = ~n_223 & ~n_276;
assign n_278 = ~n_275 &  n_277;
assign n_279 = ~n_223 & ~n_278;
assign n_280 = ~n_216 & ~n_218;
assign n_281 = ~n_219 & ~n_280;
assign n_282 = ~n_279 &  n_281;
assign n_283 = ~n_219 & ~n_282;
assign n_284 = ~n_6 &  n_214;
assign n_285 = ~n_215 & ~n_284;
assign n_286 = ~n_283 &  n_285;
assign n_287 = ~n_215 & ~n_286;
assign n_288 =  n_5 & ~n_287;
assign n_289 =  i2[11] &  i1[14];
assign n_290 =  n_283 & ~n_285;
assign n_291 = ~n_286 & ~n_290;
assign n_292 =  n_289 &  n_291;
assign n_293 =  i2[12] &  i1[14];
assign n_294 =  n_279 & ~n_281;
assign n_295 = ~n_282 & ~n_294;
assign n_296 =  n_293 &  n_295;
assign n_297 =  i2[13] &  i1[14];
assign n_298 =  n_275 & ~n_277;
assign n_299 = ~n_278 & ~n_298;
assign n_300 =  n_297 &  n_299;
assign n_301 =  i2[14] &  i1[14];
assign n_302 =  n_271 & ~n_273;
assign n_303 = ~n_274 & ~n_302;
assign n_304 =  n_301 &  n_303;
assign n_305 =  n_267 & ~n_269;
assign n_306 = ~n_270 & ~n_305;
assign n_307 =  i2[15] &  i1[14];
assign n_308 =  n_306 &  n_307;
assign n_309 =  n_263 & ~n_265;
assign n_310 = ~n_266 & ~n_309;
assign n_311 =  i2[16] &  i1[14];
assign n_312 =  n_310 &  n_311;
assign n_313 =  n_259 & ~n_261;
assign n_314 = ~n_262 & ~n_313;
assign n_315 =  i2[17] &  i1[14];
assign n_316 =  n_314 &  n_315;
assign n_317 =  n_255 & ~n_257;
assign n_318 = ~n_258 & ~n_317;
assign n_319 =  i2[18] &  i1[14];
assign n_320 =  n_318 &  n_319;
assign n_321 = ~n_251 & ~n_253;
assign n_322 = ~n_254 & ~n_321;
assign n_323 =  i2[19] &  i1[14];
assign n_324 =  n_322 &  n_323;
assign n_325 = ~n_318 & ~n_319;
assign n_326 = ~n_320 & ~n_325;
assign n_327 =  n_324 &  n_326;
assign n_328 = ~n_320 & ~n_327;
assign n_329 = ~n_314 & ~n_315;
assign n_330 = ~n_316 & ~n_329;
assign n_331 = ~n_328 &  n_330;
assign n_332 = ~n_316 & ~n_331;
assign n_333 = ~n_310 & ~n_311;
assign n_334 = ~n_312 & ~n_333;
assign n_335 = ~n_332 &  n_334;
assign n_336 = ~n_312 & ~n_335;
assign n_337 = ~n_306 & ~n_307;
assign n_338 = ~n_308 & ~n_337;
assign n_339 = ~n_336 &  n_338;
assign n_340 = ~n_308 & ~n_339;
assign n_341 = ~n_301 & ~n_303;
assign n_342 = ~n_304 & ~n_341;
assign n_343 = ~n_340 &  n_342;
assign n_344 = ~n_304 & ~n_343;
assign n_345 = ~n_297 & ~n_299;
assign n_346 = ~n_300 & ~n_345;
assign n_347 = ~n_344 &  n_346;
assign n_348 = ~n_300 & ~n_347;
assign n_349 = ~n_293 & ~n_295;
assign n_350 = ~n_296 & ~n_349;
assign n_351 = ~n_348 &  n_350;
assign n_352 = ~n_296 & ~n_351;
assign n_353 = ~n_289 & ~n_291;
assign n_354 = ~n_292 & ~n_353;
assign n_355 = ~n_352 &  n_354;
assign n_356 = ~n_292 & ~n_355;
assign n_357 = ~n_5 &  n_287;
assign n_358 = ~n_288 & ~n_357;
assign n_359 = ~n_356 &  n_358;
assign n_360 = ~n_288 & ~n_359;
assign n_361 =  n_4 & ~n_360;
assign n_362 =  i2[11] &  i1[13];
assign n_363 =  n_356 & ~n_358;
assign n_364 = ~n_359 & ~n_363;
assign n_365 =  n_362 &  n_364;
assign n_366 =  i2[12] &  i1[13];
assign n_367 =  n_352 & ~n_354;
assign n_368 = ~n_355 & ~n_367;
assign n_369 =  n_366 &  n_368;
assign n_370 =  i2[13] &  i1[13];
assign n_371 =  n_348 & ~n_350;
assign n_372 = ~n_351 & ~n_371;
assign n_373 =  n_370 &  n_372;
assign n_374 =  i2[14] &  i1[13];
assign n_375 =  n_344 & ~n_346;
assign n_376 = ~n_347 & ~n_375;
assign n_377 =  n_374 &  n_376;
assign n_378 =  i2[15] &  i1[13];
assign n_379 =  n_340 & ~n_342;
assign n_380 = ~n_343 & ~n_379;
assign n_381 =  n_378 &  n_380;
assign n_382 =  n_336 & ~n_338;
assign n_383 = ~n_339 & ~n_382;
assign n_384 =  i2[16] &  i1[13];
assign n_385 =  n_383 &  n_384;
assign n_386 =  n_332 & ~n_334;
assign n_387 = ~n_335 & ~n_386;
assign n_388 =  i2[17] &  i1[13];
assign n_389 =  n_387 &  n_388;
assign n_390 =  n_328 & ~n_330;
assign n_391 = ~n_331 & ~n_390;
assign n_392 =  i2[18] &  i1[13];
assign n_393 =  n_391 &  n_392;
assign n_394 = ~n_324 & ~n_326;
assign n_395 = ~n_327 & ~n_394;
assign n_396 =  i2[19] &  i1[13];
assign n_397 =  n_395 &  n_396;
assign n_398 = ~n_391 & ~n_392;
assign n_399 = ~n_393 & ~n_398;
assign n_400 =  n_397 &  n_399;
assign n_401 = ~n_393 & ~n_400;
assign n_402 = ~n_387 & ~n_388;
assign n_403 = ~n_389 & ~n_402;
assign n_404 = ~n_401 &  n_403;
assign n_405 = ~n_389 & ~n_404;
assign n_406 = ~n_383 & ~n_384;
assign n_407 = ~n_385 & ~n_406;
assign n_408 = ~n_405 &  n_407;
assign n_409 = ~n_385 & ~n_408;
assign n_410 = ~n_378 & ~n_380;
assign n_411 = ~n_381 & ~n_410;
assign n_412 = ~n_409 &  n_411;
assign n_413 = ~n_381 & ~n_412;
assign n_414 = ~n_374 & ~n_376;
assign n_415 = ~n_377 & ~n_414;
assign n_416 = ~n_413 &  n_415;
assign n_417 = ~n_377 & ~n_416;
assign n_418 = ~n_370 & ~n_372;
assign n_419 = ~n_373 & ~n_418;
assign n_420 = ~n_417 &  n_419;
assign n_421 = ~n_373 & ~n_420;
assign n_422 = ~n_366 & ~n_368;
assign n_423 = ~n_369 & ~n_422;
assign n_424 = ~n_421 &  n_423;
assign n_425 = ~n_369 & ~n_424;
assign n_426 = ~n_362 & ~n_364;
assign n_427 = ~n_365 & ~n_426;
assign n_428 = ~n_425 &  n_427;
assign n_429 = ~n_365 & ~n_428;
assign n_430 = ~n_4 &  n_360;
assign n_431 = ~n_361 & ~n_430;
assign n_432 = ~n_429 &  n_431;
assign n_433 = ~n_361 & ~n_432;
assign n_434 =  n_3 & ~n_433;
assign n_435 =  i2[11] &  i1[12];
assign n_436 =  n_429 & ~n_431;
assign n_437 = ~n_432 & ~n_436;
assign n_438 =  n_435 &  n_437;
assign n_439 =  i2[12] &  i1[12];
assign n_440 =  n_425 & ~n_427;
assign n_441 = ~n_428 & ~n_440;
assign n_442 =  n_439 &  n_441;
assign n_443 =  i2[13] &  i1[12];
assign n_444 =  n_421 & ~n_423;
assign n_445 = ~n_424 & ~n_444;
assign n_446 =  n_443 &  n_445;
assign n_447 =  i2[14] &  i1[12];
assign n_448 =  n_417 & ~n_419;
assign n_449 = ~n_420 & ~n_448;
assign n_450 =  n_447 &  n_449;
assign n_451 =  i2[15] &  i1[12];
assign n_452 =  n_413 & ~n_415;
assign n_453 = ~n_416 & ~n_452;
assign n_454 =  n_451 &  n_453;
assign n_455 =  i2[16] &  i1[12];
assign n_456 =  n_409 & ~n_411;
assign n_457 = ~n_412 & ~n_456;
assign n_458 =  n_455 &  n_457;
assign n_459 =  n_405 & ~n_407;
assign n_460 = ~n_408 & ~n_459;
assign n_461 =  i2[17] &  i1[12];
assign n_462 =  n_460 &  n_461;
assign n_463 =  n_401 & ~n_403;
assign n_464 = ~n_404 & ~n_463;
assign n_465 =  i2[18] &  i1[12];
assign n_466 =  n_464 &  n_465;
assign n_467 = ~n_397 & ~n_399;
assign n_468 = ~n_400 & ~n_467;
assign n_469 =  i2[19] &  i1[12];
assign n_470 =  n_468 &  n_469;
assign n_471 = ~n_464 & ~n_465;
assign n_472 = ~n_466 & ~n_471;
assign n_473 =  n_470 &  n_472;
assign n_474 = ~n_466 & ~n_473;
assign n_475 = ~n_460 & ~n_461;
assign n_476 = ~n_462 & ~n_475;
assign n_477 = ~n_474 &  n_476;
assign n_478 = ~n_462 & ~n_477;
assign n_479 = ~n_455 & ~n_457;
assign n_480 = ~n_458 & ~n_479;
assign n_481 = ~n_478 &  n_480;
assign n_482 = ~n_458 & ~n_481;
assign n_483 = ~n_451 & ~n_453;
assign n_484 = ~n_454 & ~n_483;
assign n_485 = ~n_482 &  n_484;
assign n_486 = ~n_454 & ~n_485;
assign n_487 = ~n_447 & ~n_449;
assign n_488 = ~n_450 & ~n_487;
assign n_489 = ~n_486 &  n_488;
assign n_490 = ~n_450 & ~n_489;
assign n_491 = ~n_443 & ~n_445;
assign n_492 = ~n_446 & ~n_491;
assign n_493 = ~n_490 &  n_492;
assign n_494 = ~n_446 & ~n_493;
assign n_495 = ~n_439 & ~n_441;
assign n_496 = ~n_442 & ~n_495;
assign n_497 = ~n_494 &  n_496;
assign n_498 = ~n_442 & ~n_497;
assign n_499 = ~n_435 & ~n_437;
assign n_500 = ~n_438 & ~n_499;
assign n_501 = ~n_498 &  n_500;
assign n_502 = ~n_438 & ~n_501;
assign n_503 = ~n_3 &  n_433;
assign n_504 = ~n_434 & ~n_503;
assign n_505 = ~n_502 &  n_504;
assign n_506 = ~n_434 & ~n_505;
assign n_507 =  n_2 & ~n_506;
assign n_508 =  i2[11] &  i1[11];
assign n_509 =  n_502 & ~n_504;
assign n_510 = ~n_505 & ~n_509;
assign n_511 =  n_508 &  n_510;
assign n_512 =  i2[12] &  i1[11];
assign n_513 =  n_498 & ~n_500;
assign n_514 = ~n_501 & ~n_513;
assign n_515 =  n_512 &  n_514;
assign n_516 =  i2[13] &  i1[11];
assign n_517 =  n_494 & ~n_496;
assign n_518 = ~n_497 & ~n_517;
assign n_519 =  n_516 &  n_518;
assign n_520 =  i2[14] &  i1[11];
assign n_521 =  n_490 & ~n_492;
assign n_522 = ~n_493 & ~n_521;
assign n_523 =  n_520 &  n_522;
assign n_524 =  i2[15] &  i1[11];
assign n_525 =  n_486 & ~n_488;
assign n_526 = ~n_489 & ~n_525;
assign n_527 =  n_524 &  n_526;
assign n_528 =  i2[16] &  i1[11];
assign n_529 =  n_482 & ~n_484;
assign n_530 = ~n_485 & ~n_529;
assign n_531 =  n_528 &  n_530;
assign n_532 =  i2[17] &  i1[11];
assign n_533 =  n_478 & ~n_480;
assign n_534 = ~n_481 & ~n_533;
assign n_535 =  n_532 &  n_534;
assign n_536 =  n_474 & ~n_476;
assign n_537 = ~n_477 & ~n_536;
assign n_538 =  i2[18] &  i1[11];
assign n_539 =  n_537 &  n_538;
assign n_540 = ~n_470 & ~n_472;
assign n_541 = ~n_473 & ~n_540;
assign n_542 =  i2[19] &  i1[11];
assign n_543 =  n_541 &  n_542;
assign n_544 = ~n_537 & ~n_538;
assign n_545 = ~n_539 & ~n_544;
assign n_546 =  n_543 &  n_545;
assign n_547 = ~n_539 & ~n_546;
assign n_548 = ~n_532 & ~n_534;
assign n_549 = ~n_535 & ~n_548;
assign n_550 = ~n_547 &  n_549;
assign n_551 = ~n_535 & ~n_550;
assign n_552 = ~n_528 & ~n_530;
assign n_553 = ~n_531 & ~n_552;
assign n_554 = ~n_551 &  n_553;
assign n_555 = ~n_531 & ~n_554;
assign n_556 = ~n_524 & ~n_526;
assign n_557 = ~n_527 & ~n_556;
assign n_558 = ~n_555 &  n_557;
assign n_559 = ~n_527 & ~n_558;
assign n_560 = ~n_520 & ~n_522;
assign n_561 = ~n_523 & ~n_560;
assign n_562 = ~n_559 &  n_561;
assign n_563 = ~n_523 & ~n_562;
assign n_564 = ~n_516 & ~n_518;
assign n_565 = ~n_519 & ~n_564;
assign n_566 = ~n_563 &  n_565;
assign n_567 = ~n_519 & ~n_566;
assign n_568 = ~n_512 & ~n_514;
assign n_569 = ~n_515 & ~n_568;
assign n_570 = ~n_567 &  n_569;
assign n_571 = ~n_515 & ~n_570;
assign n_572 = ~n_508 & ~n_510;
assign n_573 = ~n_511 & ~n_572;
assign n_574 = ~n_571 &  n_573;
assign n_575 = ~n_511 & ~n_574;
assign n_576 = ~n_2 &  n_506;
assign n_577 = ~n_507 & ~n_576;
assign n_578 = ~n_575 &  n_577;
assign n_579 = ~n_507 & ~n_578;
assign n_580 =  n_1 & ~n_579;
assign n_581 =  i2[11] &  i1[10];
assign n_582 =  n_575 & ~n_577;
assign n_583 = ~n_578 & ~n_582;
assign n_584 =  n_581 &  n_583;
assign n_585 =  i2[12] &  i1[10];
assign n_586 =  n_571 & ~n_573;
assign n_587 = ~n_574 & ~n_586;
assign n_588 =  n_585 &  n_587;
assign n_589 =  i2[13] &  i1[10];
assign n_590 =  n_567 & ~n_569;
assign n_591 = ~n_570 & ~n_590;
assign n_592 =  n_589 &  n_591;
assign n_593 =  i2[14] &  i1[10];
assign n_594 =  n_563 & ~n_565;
assign n_595 = ~n_566 & ~n_594;
assign n_596 =  n_593 &  n_595;
assign n_597 =  i2[15] &  i1[10];
assign n_598 =  n_559 & ~n_561;
assign n_599 = ~n_562 & ~n_598;
assign n_600 =  n_597 &  n_599;
assign n_601 =  i2[16] &  i1[10];
assign n_602 =  n_555 & ~n_557;
assign n_603 = ~n_558 & ~n_602;
assign n_604 =  n_601 &  n_603;
assign n_605 =  i2[17] &  i1[10];
assign n_606 =  n_551 & ~n_553;
assign n_607 = ~n_554 & ~n_606;
assign n_608 =  n_605 &  n_607;
assign n_609 =  i2[18] &  i1[10];
assign n_610 =  n_547 & ~n_549;
assign n_611 = ~n_550 & ~n_610;
assign n_612 =  n_609 &  n_611;
assign n_613 = ~n_543 & ~n_545;
assign n_614 = ~n_546 & ~n_613;
assign n_615 =  i2[19] &  i1[10];
assign n_616 =  n_614 &  n_615;
assign n_617 = ~n_609 & ~n_611;
assign n_618 = ~n_612 & ~n_617;
assign n_619 =  n_616 &  n_618;
assign n_620 = ~n_612 & ~n_619;
assign n_621 = ~n_605 & ~n_607;
assign n_622 = ~n_608 & ~n_621;
assign n_623 = ~n_620 &  n_622;
assign n_624 = ~n_608 & ~n_623;
assign n_625 = ~n_601 & ~n_603;
assign n_626 = ~n_604 & ~n_625;
assign n_627 = ~n_624 &  n_626;
assign n_628 = ~n_604 & ~n_627;
assign n_629 = ~n_597 & ~n_599;
assign n_630 = ~n_600 & ~n_629;
assign n_631 = ~n_628 &  n_630;
assign n_632 = ~n_600 & ~n_631;
assign n_633 = ~n_593 & ~n_595;
assign n_634 = ~n_596 & ~n_633;
assign n_635 = ~n_632 &  n_634;
assign n_636 = ~n_596 & ~n_635;
assign n_637 = ~n_589 & ~n_591;
assign n_638 = ~n_592 & ~n_637;
assign n_639 = ~n_636 &  n_638;
assign n_640 = ~n_592 & ~n_639;
assign n_641 = ~n_585 & ~n_587;
assign n_642 = ~n_588 & ~n_641;
assign n_643 = ~n_640 &  n_642;
assign n_644 = ~n_588 & ~n_643;
assign n_645 = ~n_581 & ~n_583;
assign n_646 = ~n_584 & ~n_645;
assign n_647 = ~n_644 &  n_646;
assign n_648 = ~n_584 & ~n_647;
assign n_649 = ~n_1 &  n_579;
assign n_650 = ~n_580 & ~n_649;
assign n_651 = ~n_648 &  n_650;
assign n_652 = ~n_580 & ~n_651;
assign n_653 =  a[0] &  n_652;
assign n_654 = ~a[0] & ~n_652;
assign n_655 =  n_648 & ~n_650;
assign n_656 = ~n_651 & ~n_655;
assign n_657 = ~a[1] &  n_656;
assign n_658 =  a[1] & ~n_656;
assign n_659 =  n_644 & ~n_646;
assign n_660 = ~n_647 & ~n_659;
assign n_661 = ~a[2] &  n_660;
assign n_662 =  a[2] & ~n_660;
assign n_663 =  n_640 & ~n_642;
assign n_664 = ~n_643 & ~n_663;
assign n_665 = ~a[3] &  n_664;
assign n_666 =  a[3] & ~n_664;
assign n_667 =  n_636 & ~n_638;
assign n_668 = ~n_639 & ~n_667;
assign n_669 = ~a[4] &  n_668;
assign n_670 =  a[4] & ~n_668;
assign n_671 =  n_632 & ~n_634;
assign n_672 = ~n_635 & ~n_671;
assign n_673 = ~a[5] &  n_672;
assign n_674 =  a[5] & ~n_672;
assign n_675 =  n_628 & ~n_630;
assign n_676 = ~n_631 & ~n_675;
assign n_677 = ~a[6] &  n_676;
assign n_678 =  a[6] & ~n_676;
assign n_679 =  n_624 & ~n_626;
assign n_680 = ~n_627 & ~n_679;
assign n_681 = ~a[7] &  n_680;
assign n_682 =  a[7] & ~n_680;
assign n_683 =  n_620 & ~n_622;
assign n_684 = ~n_623 & ~n_683;
assign n_685 = ~a[8] &  n_684;
assign n_686 =  a[8] & ~n_684;
assign n_687 = ~n_616 & ~n_618;
assign n_688 = ~n_619 & ~n_687;
assign n_689 = ~a[9] &  n_688;
assign n_690 =  a[9] & ~n_688;
assign n_691 = ~n_614 & ~n_615;
assign n_692 = ~n_616 & ~n_691;
assign n_693 = ~a[10] &  n_692;
assign n_694 =  a[10] & ~n_692;
assign n_695 = ~n_541 & ~n_542;
assign n_696 = ~n_543 & ~n_695;
assign n_697 = ~a[11] &  n_696;
assign n_698 =  a[11] & ~n_696;
assign n_699 = ~n_468 & ~n_469;
assign n_700 = ~n_470 & ~n_699;
assign n_701 = ~a[12] &  n_700;
assign n_702 =  a[12] & ~n_700;
assign n_703 = ~n_395 & ~n_396;
assign n_704 = ~n_397 & ~n_703;
assign n_705 = ~a[13] &  n_704;
assign n_706 =  a[13] & ~n_704;
assign n_707 = ~n_322 & ~n_323;
assign n_708 = ~n_324 & ~n_707;
assign n_709 = ~a[14] &  n_708;
assign n_710 =  a[14] & ~n_708;
assign n_711 = ~n_249 & ~n_250;
assign n_712 = ~n_251 & ~n_711;
assign n_713 = ~a[15] &  n_712;
assign n_714 =  a[15] & ~n_712;
assign n_715 = ~n_176 & ~n_177;
assign n_716 = ~n_178 & ~n_715;
assign n_717 = ~a[16] &  n_716;
assign n_718 =  a[16] & ~n_716;
assign n_719 = ~n_100 & ~n_104;
assign n_720 = ~n_105 & ~n_719;
assign n_721 = ~a[17] &  n_720;
assign n_722 =  a[17] & ~n_720;
assign n_723 = ~n_30 & ~n_31;
assign n_724 = ~n_32 & ~n_723;
assign n_725 = ~a[18] &  n_724;
assign n_726 =  i2[19] &  i1[19];
assign n_727 = ~a[19] & ~n_726;
assign n_728 =  a[19] &  n_726;
assign n_729 = ~n_727 & ~n_728;
assign n_730 =  a[18] & ~n_724;
assign n_731 = ~n_729 & ~n_730;
assign n_732 = ~n_725 &  n_731;
assign n_733 = ~i1[15] & ~i1[14];
assign n_734 = ~i1[13] & ~i1[12];
assign n_735 =  n_733 &  n_734;
assign n_736 =  i1[19] & ~i1[18];
assign n_737 = ~i1[17] & ~i1[16];
assign n_738 =  n_736 &  n_737;
assign n_739 =  n_735 &  n_738;
assign n_740 = ~i1[11] & ~i1[10];
assign n_741 =  n_739 &  n_740;
assign n_742 = ~i2[15] & ~i2[14];
assign n_743 = ~i2[13] & ~i2[12];
assign n_744 =  n_742 &  n_743;
assign n_745 =  i2[19] & ~i2[18];
assign n_746 = ~i2[17] & ~i2[16];
assign n_747 =  n_745 &  n_746;
assign n_748 =  n_744 &  n_747;
assign n_749 = ~i2[11] & ~i2[10];
assign n_750 =  n_748 &  n_749;
assign n_751 = ~n_741 & ~n_750;
assign n_752 =  n_732 &  n_751;
assign n_753 = ~n_722 &  n_752;
assign n_754 = ~n_721 &  n_753;
assign n_755 = ~n_718 &  n_754;
assign n_756 = ~n_717 &  n_755;
assign n_757 = ~n_714 &  n_756;
assign n_758 = ~n_713 &  n_757;
assign n_759 = ~n_710 &  n_758;
assign n_760 = ~n_709 &  n_759;
assign n_761 = ~n_706 &  n_760;
assign n_762 = ~n_705 &  n_761;
assign n_763 = ~n_702 &  n_762;
assign n_764 = ~n_701 &  n_763;
assign n_765 = ~n_698 &  n_764;
assign n_766 = ~n_697 &  n_765;
assign n_767 = ~n_694 &  n_766;
assign n_768 = ~n_693 &  n_767;
assign n_769 = ~n_690 &  n_768;
assign n_770 = ~n_689 &  n_769;
assign n_771 = ~n_686 &  n_770;
assign n_772 = ~n_685 &  n_771;
assign n_773 = ~n_682 &  n_772;
assign n_774 = ~n_681 &  n_773;
assign n_775 = ~n_678 &  n_774;
assign n_776 = ~n_677 &  n_775;
assign n_777 = ~n_674 &  n_776;
assign n_778 = ~n_673 &  n_777;
assign n_779 = ~n_670 &  n_778;
assign n_780 = ~n_669 &  n_779;
assign n_781 = ~n_666 &  n_780;
assign n_782 = ~n_665 &  n_781;
assign n_783 = ~n_662 &  n_782;
assign n_784 = ~n_661 &  n_783;
assign n_785 = ~n_658 &  n_784;
assign n_786 = ~n_657 &  n_785;
assign n_787 = ~n_654 &  n_786;
assign n_788 = ~n_653 &  n_787;
assign o_1 =  n_788;
endmodule

