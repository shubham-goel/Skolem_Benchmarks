// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module neclaftp3002_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, x_181, x_182, x_183, x_184, x_185, x_186, x_187, x_188, x_189, x_190, x_191, x_192, x_193, x_194, x_195, x_196, x_197, x_198, x_199, x_200, x_201, x_202, x_203, x_204, x_205, x_206, x_207, x_208, x_209, x_210, x_211, x_212, x_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, x_460, x_461, x_462, x_463, x_464, x_465, x_466, x_467, x_468, x_469, x_470, x_471, x_472, x_473, x_474, x_475, x_476, x_477, x_478, x_479, x_480, x_481, x_482, x_483, x_484, x_485, x_486, x_487, x_488, x_489, x_490, x_491, x_492, x_493, x_494, x_495, x_496, x_497, x_498, x_499, x_500, x_501, x_502, x_503, x_504, x_505, x_506, x_507, x_508, x_509, x_510, x_511, x_512, x_513, x_514, x_515, x_516, x_517, x_518, x_519, x_520, x_521, x_522, x_523, x_524, x_525, x_526, x_527, x_528, x_529, x_530, x_531, x_532, x_533, x_534, x_535, x_536, x_537, x_538, x_539, x_540, x_541, x_542, x_543, x_544, x_545, x_546, x_547, x_548, x_549, x_550, x_551, x_552, x_553, x_554, x_555, x_556, x_557, x_558, x_559, x_560, x_561, x_562, x_563, x_564, x_565, x_566, x_567, x_568, x_569, x_570, x_571, x_572, x_573, x_574, x_575, x_576, x_577, x_578, x_579, x_580, x_581, x_582, x_583, x_584, x_585, x_586, x_587, x_588, x_589, x_590, x_591, x_592, x_593, x_594, x_595, x_596, x_597, x_598, x_599, x_600, x_601, x_602, x_603, x_604, x_605, x_606, x_607, x_608, x_609, x_610, x_611, x_612, x_613, x_614, x_615, x_616, x_617, x_618, x_619, x_620, x_621, x_622, x_623, x_624, x_625, x_626, x_627, x_628, x_629, x_630, x_631, x_632, x_633, x_634, x_635, x_636, x_637, x_638, x_639, x_640, x_641, x_642, x_643, x_644, x_645, x_646, x_647, x_648, x_649, x_650, x_651, x_652, x_653, x_654, x_655, x_656, x_657, x_658, x_659, x_660, x_661, x_662, x_663, x_664, x_665, x_666, x_667, x_668, x_669, x_670, x_671, x_672, x_673, x_674, x_675, x_676, x_677, x_678, x_679, x_680, x_681, x_682, x_683, x_684, x_685, x_686, x_687, x_688, x_689, x_690, x_691, x_692, x_693, x_694, x_695, x_696, x_697, x_698, x_699, x_700, x_701, x_702, x_703, x_704, x_705, x_706, x_707, x_708, x_709, x_710, x_711, x_712, x_713, x_714, x_715, x_716, x_717, x_718, x_719, x_720, x_721, x_722, x_723, x_724, x_725, x_726, x_727, x_728, x_729, x_730, x_731, x_732, x_733, x_734, x_735, x_736, x_737, x_738, x_739, x_740, x_741, x_742, x_743, x_744, x_745, x_746, x_747, x_748, x_749, x_750, x_751, x_752, x_753, x_754, x_755, x_756, x_757, x_758, x_759, x_760, x_761, x_762, x_763, x_764, x_765, x_766, x_767, x_768, x_769, x_770, x_771, x_772, x_773, x_774, x_775, x_776, x_777, x_778, x_779, x_780, x_781, x_782, x_783, x_784, x_785, x_786, x_787, x_788, x_789, x_790, x_791, x_792, x_793, x_794, x_795, x_796, x_797, x_798, x_799, x_800, x_801, x_802, x_803, x_804, x_805, x_806, x_807, x_808, x_809, x_810, x_811, x_812, x_813, x_814, x_815, x_816, x_817, x_818, x_819, x_820, x_821, x_822, x_823, x_824, x_825, x_826, x_827, x_828, x_829, x_830, x_831, x_832, x_833, x_834, x_835, x_836, x_837, x_838, x_839, x_840, x_841, x_842, x_843, x_844, x_845, x_846, x_847, x_848, x_849, x_850, x_851, x_852, x_853, x_854, x_855, x_856, x_857, x_858, x_859, x_860, x_861, x_862, x_863, x_864, x_865, x_866, x_867, x_868, x_869, x_870, x_871, x_872, x_873, x_874, x_875, x_876, x_877, x_878, x_879, x_880, x_881, x_882, x_883, x_884, x_885, x_886, x_887, x_888, x_889, x_890, x_891, x_892, x_893, x_894, x_895, x_896, x_897, x_898, x_899, x_900, x_901, x_902, x_903, x_904, x_905, x_906, x_907, x_908, x_909, x_910, x_911, x_912, x_913, x_914, x_915, x_916, x_917, x_918, x_919, x_920, x_921, x_922, x_923, x_924, x_925, x_926, x_927, x_928, x_929, x_930, x_931, x_932, x_933, x_934, x_935, x_936, x_937, x_938, x_939, x_940, x_941, x_942, x_943, x_944, x_945, x_946, x_947, x_948, x_949, x_950, x_951, x_952, x_953, x_954, x_955, x_956, x_957, x_958, x_959, x_960, x_961, x_962, x_963, x_964, x_965, x_966, x_967, x_968, x_969, x_970, x_971, x_972, x_973, x_974, x_975, x_976, x_977, x_978, x_979, x_980, x_981, x_982, x_983, x_984, x_985, x_986, x_987, x_988, x_989, x_990, x_991, x_992, x_993, x_994, x_995, x_996, x_997, x_998, x_999, x_1000, x_1001, x_1002, x_1003, x_1004, x_1005, x_1006, x_1007, x_1008, x_1009, x_1010, x_1011, x_1012, x_1013, x_1014, x_1015, x_1016, x_1017, x_1018, x_1019, x_1020, x_1021, x_1022, x_1023, x_1024, x_1025, x_1026, x_1027, x_1028, x_1029, x_1030, x_1031, x_1032, x_1033, x_1034, x_1035, x_1036, x_1037, x_1038, x_1039, x_1040, x_1041, x_1042, x_1043, x_1044, x_1045, x_1046, x_1047, x_1048, x_1049, x_1050, x_1051, x_1052, x_1053, x_1054, x_1055, x_1056, x_1057, x_1058, x_1059, x_1060, x_1061, x_1062, x_1063, x_1064, x_1065, x_1066, x_1067, x_1068, x_1069, x_1070, x_1071, x_1072, x_1073, x_1074, x_1075, x_1076, x_1077, x_1078, x_1079, x_1080, x_1081, x_1082, x_1083, x_1084, x_1085, x_1086, x_1087, x_1088, x_1089, x_1090, x_1091, x_1092, x_1093, x_1094, x_1095, x_1096, x_1097, x_1098, x_1099, x_1100, x_1101, x_1102, x_1103, x_1104, x_1105, x_1106, x_1107, x_1108, x_1109, x_1110, x_1111, x_1112, x_1113, x_1114, x_1115, x_1116, x_1117, x_1118, x_1119, x_1120, x_1121, x_1122, x_1123, x_1124, x_1125, x_1126, x_1127, x_1128, x_1129, x_1130, x_1131, x_1132, x_1133, x_1134, x_1135, x_1136, x_1137, x_1138, x_1139, x_1140, x_1141, x_1142, x_1143, x_1144, x_1145, x_1146, x_1147, x_1148, x_1149, x_1150, x_1151, x_1152, x_1153, x_1154, x_1155, x_1156, x_1157, x_1158, x_1159, x_1160, x_1161, x_1162, x_1163, x_1164, x_1165, x_1166, x_1167, x_1168, x_1169, x_1170, x_1171, x_1172, x_1173, x_1174, x_1175, x_1176, x_1177, x_1178, x_1179, x_1180, x_1181, x_1182, x_1183, x_1184, x_1185, x_1186, x_1187, x_1188, x_1189, x_1190, x_1191, x_1192, x_1193, x_1194, x_1195, x_1196, x_1197, x_1198, x_1199, x_1200, x_1201, x_1202, x_1203, x_1204, x_1205, x_1206, x_1207, x_1208, x_1209, x_1210, x_1211, x_1212, x_1213, x_1214, x_1215, x_1216, x_1217, x_1218, x_1219, x_1220, x_1221, x_1222, x_1223, x_1224, x_1225, x_1226, x_1227, x_1228, x_1229, x_1230, x_1231, x_1232, x_1233, x_1234, x_1235, x_1236, x_1237, x_1238, x_1239, x_1240, x_1241, x_1242, x_1243, x_1244, x_1245, x_1246, x_1247, x_1248, x_1249, x_1250, x_1251, x_1252, x_1253, x_1254, x_1255, x_1256, x_1257, x_1258, x_1259, x_1260, x_1261, x_1262, x_1263, x_1264, x_1265, x_1266, x_1267, x_1268, x_1269, x_1270, x_1271, x_1272, x_1273, x_1274, x_1275, x_1276, x_1277, x_1278, x_1279, x_1280, x_1281, x_1282, x_1283, x_1284, x_1285, x_1286, x_1287, x_1288, x_1289, x_1290, x_1291, x_1292, x_1293, x_1294, x_1295, x_1296, x_1297, x_1298, x_1299, x_1300, x_1301, x_1302, x_1303, x_1304, x_1305, x_1306, x_1307, x_1308, x_1309, x_1310, x_1311, x_1312, x_1313, x_1314, x_1315, x_1316, x_1317, x_1318, x_1319, x_1320, x_1321, x_1322, x_1323, x_1324, x_1325, x_1326, x_1327, x_1328, x_1329, x_1330, x_1331, x_1332, x_1333, x_1334, x_1335, x_1336, x_1337, x_1338, x_1339, x_1340, x_1341, x_1342, x_1343, x_1344, x_1345, x_1346, x_1347, x_1348, x_1349, x_1350, x_1351, x_1352, x_1353, x_1354, x_1355, x_1356, x_1357, x_1358, x_1359, x_1360, x_1361, x_1362, x_1363, x_1364, x_1365, x_1366, x_1367, x_1368, x_1369, x_1370, x_1371, x_1372, x_1373, x_1374, x_1375, x_1376, x_1377, x_1378, x_1379, x_1380, x_1381, x_1382, x_1383, x_1384, x_1385, x_1386, x_1387, x_1388, x_1389, x_1390, x_1391, x_1392, x_1393, x_1394, x_1395, x_1396, x_1397, x_1398, x_1399, x_1400, x_1401, x_1402, x_1403, x_1404, x_1405, x_1406, x_1407, x_1408, x_1409, x_1410, x_1411, x_1412, x_1413, x_1414, x_1415, x_1416, x_1417, x_1418, x_1419, x_1420, x_1421, x_1422, x_1423, x_1424, x_1425, x_1426, x_1427, x_1428, x_1429, x_1430, x_1431, x_1432, x_1433, x_1434, x_1435, x_1436, x_1437, x_1438, x_1439, x_1440, x_1441, x_1442, x_1443, x_1444, x_1445, x_1446, x_1447, x_1448, x_1449, x_1450, x_1451, x_1452, x_1453, x_1454, x_1455, x_1456, x_1457, x_1458, x_1459, x_1460, x_1461, x_1462, x_1463, x_1464, x_1465, x_1466, x_1467, x_1468, x_1469, x_1470, x_1471, x_1472, x_1473, x_1474, x_1475, x_1476, x_1477, x_1478, x_1479, x_1480, x_1481, x_1482, x_1483, x_1484, x_1485, x_1486, x_1487, x_1488, x_1489, x_1490, x_1491, x_1492, x_1493, x_1494, x_1495, x_1496, x_1497, x_1498, x_1499, x_1500, x_1501, x_1502, x_1503, x_1504, x_1505, x_1506, x_1507, x_1508, x_1509, x_1510, x_1511, x_1512, x_1513, x_1514, x_1515, x_1516, x_1517, x_1518, x_1519, x_1520, x_1521, x_1522, x_1523, x_1524, x_1525, x_1526, x_1527, x_1528, x_1529, x_1530, x_1531, x_1532, x_1533, x_1534, x_1535, x_1536, x_1537, x_1538, x_1539, x_1540, x_1541, x_1542, x_1543, x_1544, x_1545, x_1546, x_1547, x_1548, x_1549, x_1550, x_1551, x_1552, x_1553, x_1554, x_1555, x_1556, x_1557, x_1558, x_1559, x_1560, x_1561, x_1562, x_1563, x_1564, x_1565, x_1566, x_1567, x_1568, x_1569, x_1570, x_1571, x_1572, x_1573, x_1574, x_1575, x_1576, x_1577, x_1578, x_1579, x_1580, x_1581, x_1582, x_1583, x_1584, x_1585, x_1586, x_1587, x_1588, x_1589, x_1590, x_1591, x_1592, x_1593, x_1594, x_1595, x_1596, x_1597, x_1598, x_1599, x_1600, x_1601, x_1602, x_1603, x_1604, x_1605, x_1606, x_1607, x_1608, x_1609, x_1610, x_1611, x_1612, x_1613, x_1614, x_1615, x_1616, x_1617, x_1618, x_1619, x_1620, x_1621, x_1622, x_1623, x_1624, x_1625, x_1626, x_1627, x_1628, x_1629, x_1630, x_1631, x_1632, x_1633, x_1634, x_1635, x_1636, x_1637, x_1638, x_1639, x_1640, x_1641, x_1642, x_1643, x_1644, x_1645, x_1646, x_1647, x_1648, x_1649, x_1650, x_1651, x_1652, x_1653, x_1654, x_1655, x_1656, x_1657, x_1658, x_1659, x_1660, x_1661, x_1662, x_1663, x_1664, x_1665, x_1666, x_1667, x_1668, x_1669, x_1670, x_1671, x_1672, x_1673, x_1674, x_1675, x_1676, x_1677, x_1678, x_1679, x_1680, x_1681, x_1682, x_1683, x_1684, x_1685, x_1686, x_1687, x_1688, x_1689, x_1690, x_1691, x_1692, x_1693, x_1694, x_1695, x_1696, x_1697, x_1698, x_1699, x_1700, x_1701, x_1702, x_1703, x_1704, x_1705, x_1706, x_1707, x_1708, x_1709, x_1710, x_1711, x_1712, x_1713, x_1714, x_1715, x_1716, x_1717, x_1718, x_1719, x_1720, x_1721, x_1722, x_1723, x_1724, x_1725, x_1726, x_1727, x_1728, x_1729, x_1730, x_1731, x_1732, x_1733, x_1734, x_1735, x_1736, x_1737, x_1738, x_1739, x_1740, x_1741, x_1742, x_1743, x_1744, x_1745, x_1746, x_1747, x_1748, x_1749, x_1750, x_1751, x_1752, x_1753, x_1754, x_1755, x_1756, x_1757, x_1758, x_1759, x_1760, x_1761, x_1762, x_1763, x_1764, x_1765, x_1766, x_1767, x_1768, x_1769, x_1770, x_1771, x_1772, x_1773, x_1774, x_1775, x_1776, x_1777, x_1778, x_1779, x_1780, x_1781, x_1782, x_1783, x_1784, x_1785, x_1786, x_1787, x_1788, x_1789, x_1790, x_1791, x_1792, x_1793, x_1794, x_1795, x_1796, x_1797, x_1798, x_1799, x_1800, x_1801, x_1802, x_1803, x_1804, x_1805, x_1806, x_1807, x_1808, x_1809, x_1810, x_1811, x_1812, x_1813, x_1814, x_1815, x_1816, x_1817, x_1818, x_1819, x_1820, x_1821, x_1822, x_1823, x_1824, x_1825, x_1826, x_1827, x_1828, x_1829, x_1830, x_1831, x_1832, x_1833, x_1834, x_1835, x_1836, x_1837, x_1838, x_1839, x_1840, x_1841, x_1842, x_1843, x_1844, x_1845, x_1846, x_1847, x_1848, x_1849, x_1850, x_1851, x_1852, x_1853, x_1854, x_1855, x_1856, x_1857, x_1858, x_1859, x_1860, x_1861, x_1862, x_1863, x_1864, x_1865, x_1866, x_1867, x_1868, x_1869, x_1870, x_1871, x_1872, x_1873, x_1874, x_1875, x_1876, x_1877, x_1878, x_1879, x_1880, x_1881, x_1882, x_1883, x_1884, x_1885, x_1886, x_1887, x_1888, x_1889, x_1890, x_1891, x_1892, x_1893, x_1894, x_1895, x_1896, x_1897, x_1898, x_1899, x_1900, x_1901, x_1902, x_1903, x_1904, x_1905, x_1906, x_1907, x_1908, x_1909, x_1910, x_1911, x_1912, x_1913, x_1914, x_1915, x_1916, x_1917, x_1918, x_1919, x_1920, x_1921, x_1922, x_1923, x_1924, x_1925, x_1926, x_1927, x_1928, x_1929, x_1930, x_1931, x_1932, x_1933, x_1934, x_1935, x_1936, x_1937, x_1938, x_1939, x_1940, x_1941, x_1942, x_1943, x_1944, x_1945, x_1946, x_1947, x_1948, x_1949, x_1950, x_1951, x_1952, x_1953, x_1954, x_1955, x_1956, x_1957, x_1958, x_1959, x_1960, x_1961, x_1962, x_1963, x_1964, x_1965, x_1966, x_1967, x_1968, x_1969, x_1970, x_1971, x_1972, x_1973, x_1974, x_1975, x_1976, x_1977, x_1978, x_1979, x_1980, x_1981, x_1982, x_1983, x_1984, x_1985, x_1986, x_1987, x_1988, x_1989, x_1990, x_1991, x_1992, x_1993, x_1994, x_1995, x_1996, x_1997, x_1998, x_1999, x_2000, x_2001, x_2002, x_2003, x_2004, x_2005, x_2006, x_2007, x_2008, x_2009, x_2010, x_2011, x_2012, x_2013, x_2014, x_2015, x_2016, x_2017, x_2018, x_2019, x_2020, x_2021, x_2022, x_2023, x_2024, x_2025, x_2026, x_2027, x_2028, x_2029, x_2030, x_2031, x_2032, x_2033, x_2034, x_2035, x_2036, x_2037, x_2038, x_2039, x_2040, x_2041, x_2042, x_2043, x_2044, x_2045, x_2046, x_2047, x_2048, x_2049, x_2050, x_2051, x_2052, x_2053, x_2054, x_2055, x_2056, x_2057, x_2058, x_2059, x_2060, x_2061, x_2062, x_2063, x_2064, x_2065, x_2066, x_2067, x_2068, x_2069, x_2070, x_2071, x_2072, x_2073, x_2074, x_2075, x_2076, x_2077, x_2078, x_2079, x_2080, x_2081, x_2082, x_2083, x_2084, x_2085, x_2086, x_2087, x_2088, x_2089, x_2090, x_2091, x_2092, x_2093, x_2094, x_2095, x_2096, x_2097, x_2098, x_2099, x_2100, x_2101, x_2102, x_2103, x_2104, x_2105, x_2106, x_2107, x_2108, x_2109, x_2110, x_2111, x_2112, x_2113, x_2114, x_2115, x_2116, x_2117, x_2118, x_2119, x_2120, x_2121, x_2122, x_2123, x_2124, x_2125, x_2126, x_2127, x_2128, x_2129, x_2130, x_2131, x_2132, x_2133, x_2134, x_2135, x_2136, x_2137, x_2138, x_2139, x_2140, x_2141, x_2142, x_2143, x_2144, x_2145, x_2146, x_2147, x_2148, x_2149, x_2150, x_2151, x_2152, x_2153, x_2154, x_2155, x_2156, x_2157, x_2158, x_2159, x_2160, x_2161, x_2162, x_2163, x_2164, x_2165, x_2166, x_2167, x_2168, x_2169, x_2170, x_2171, x_2172, x_2173, x_2174, x_2175, x_2176, x_2177, x_2178, x_2179, x_2180, x_2181, x_2182, x_2183, x_2184, x_2185, x_2186, x_2187, x_2188, x_2189, x_2190, x_2191, x_2192, x_2193, x_2194, x_2195, x_2196, x_2197, x_2198, x_2199, x_2200, x_2201, x_2202, x_2203, x_2204, x_2205, x_2206, x_2207, x_2208, x_2209, x_2210, x_2211, x_2212, x_2213, x_2214, x_2215, x_2216, x_2217, x_2218, x_2219, x_2220, x_2221, x_2222, x_2223, x_2224, x_2225, x_2226, x_2227, x_2228, x_2229, x_2230, x_2231, x_2232, x_2233, x_2234, x_2235, x_2236, x_2237, x_2238, x_2239, x_2240, x_2241, x_2242, x_2243, x_2244, x_2245, x_2246, x_2247, x_2248, x_2249, x_2250, x_2251, x_2252, x_2253, x_2254, x_2255, x_2256, x_2257, x_2258, x_2259, x_2260, x_2261, x_2262, x_2263, x_2264, x_2265, x_2266, x_2267, x_2268, x_2269, x_2270, x_2271, x_2272, x_2273, x_2274, x_2275, x_2276, x_2277, x_2278, x_2279, x_2280, x_2281, x_2282, x_2283, x_2284, x_2285, x_2286, x_2287, x_2288, x_2289, x_2290, x_2291, x_2292, x_2293, x_2294, x_2295, x_2296, x_2297, x_2298, x_2299, x_2300, x_2301, x_2302, x_2303, x_2304, x_2305, x_2306, x_2307, x_2308, x_2309, x_2310, x_2311, x_2312, x_2313, x_2314, x_2315, x_2316, x_2317, x_2318, x_2319, x_2320, x_2321, x_2322, x_2323, x_2324, x_2325, x_2326, x_2327, x_2328, x_2329, x_2330, x_2331, x_2332, x_2333, x_2334, x_2335, x_2336, x_2337, x_2338, x_2339, x_2340, x_2341, x_2342, x_2343, x_2344, x_2345, x_2346, x_2347, x_2348, x_2349, x_2350, x_2351, x_2352, x_2353, x_2354, x_2355, x_2356, x_2357, x_2358, x_2359, x_2360, x_2361, x_2362, x_2363, x_2364, x_2365, x_2366, x_2367, x_2368, x_2369, x_2370, x_2371, x_2372, x_2373, x_2374, x_2375, x_2376, x_2377, x_2378, x_2379, x_2380, x_2381, x_2382, x_2383, x_2384, x_2385, x_2386, x_2387, x_2388, x_2389, x_2390, x_2391, x_2392, x_2393, x_2394, x_2395, x_2396, x_2397, x_2398, x_2399, x_2400, x_2401, x_2402, x_2403, x_2404, x_2405, x_2406, x_2407, x_2408, x_2409, x_2410, x_2411, x_2412, x_2413, x_2414, x_2415, x_2416, x_2417, x_2418, x_2419, x_2420, x_2421, x_2422, x_2423, x_2424, x_2425, x_2426, x_2427, x_2428, x_2429, x_2430, x_2431, x_2432, x_2433, x_2434, x_2435, x_2436, x_2437, x_2438, x_2439, x_2440, x_2441, x_2442, x_2443, x_2444, x_2445, x_2446, x_2447, x_2448, x_2449, x_2450, x_2451, x_2452, x_2453, x_2454, x_2455, x_2456, x_2457, x_2458, x_2459, x_2460, x_2461, x_2462, x_2463, x_2464, x_2465, x_2466, x_2467, x_2468, x_2469, x_2470, x_2471, x_2472, x_2473, x_2474, x_2475, x_2476, x_2477, x_2478, x_2479, x_2480, x_2481, x_2482, x_2483, x_2484, x_2485, x_2486, x_2487, x_2488, x_2489, x_2490, x_2491, x_2492, x_2493, x_2494, x_2495, x_2496, x_2497, x_2498, x_2499, x_2500, x_2501, x_2502, x_2503, x_2504, x_2505, x_2506, x_2507, x_2508, x_2509, x_2510, x_2511, x_2512, x_2513, x_2514, x_2515, x_2516, x_2517, x_2518, x_2519, x_2520, x_2521, x_2522, x_2523, x_2524, x_2525, x_2526, x_2527, x_2528, x_2529, x_2530, x_2531, x_2532, x_2533, x_2534, x_2535, x_2536, x_2537, x_2538, x_2539, x_2540, x_2541, x_2542, x_2543, x_2544, x_2545, x_2546, x_2547, x_2548, x_2549, x_2550, x_2551, x_2552, x_2553, x_2554, x_2555, x_2556, x_2557, x_2558, x_2559, x_2560, x_2561, x_2562, x_2563, x_2564, x_2565, x_2566, x_2567, x_2568, x_2569, x_2570, x_2571, x_2572, x_2573, x_2574, x_2575, x_2576, x_2577, x_2578, x_2579, x_2580, x_2581, x_2582, x_2583, x_2584, x_2585, x_2586, x_2587, x_2588, x_2589, x_2590, x_2591, x_2592, x_2593, x_2594, x_2595, x_2596, x_2597, x_2598, x_2599, x_2600, x_2601, x_2602, x_2603, x_2604, x_2605, x_2606, x_2607, x_2608, x_2609, x_2610, x_2611, x_2612, x_2613, x_2614, x_2615, x_2616, x_2617, x_2618, x_2619, x_2620, x_2621, x_2622, x_2623, x_2624, x_2625, x_2626, x_2627, x_2628, x_2629, x_2630, x_2631, x_2632, x_2633, x_2634, x_2635, x_2636, x_2637, x_2638, x_2639, x_2640, x_2641, x_2642, x_2643, x_2644, x_2645, x_2646, x_2647, x_2648, x_2649, x_2650, x_2651, x_2652, x_2653, x_2654, x_2655, x_2656, x_2657, x_2658, x_2659, x_2660, x_2661, x_2662, x_2663, x_2664, x_2665, x_2666, x_2667, x_2668, x_2669, x_2670, x_2671, x_2672, x_2673, x_2674, x_2675, x_2676, x_2677, x_2678, x_2679, x_2680, x_2681, x_2682, x_2683, x_2684, x_2685, x_2686, x_2687, x_2688, x_2689, x_2690, x_2691, x_2692, x_2693, x_2694, x_2695, x_2696, x_2697, x_2698, x_2699, x_2700, x_2701, x_2702, x_2703, x_2704, x_2705, x_2706, x_2707, x_2708, x_2709, x_2710, x_2711, x_2712, x_2713, x_2714, x_2715, x_2716, x_2717, x_2718, x_2719, x_2720, x_2721, x_2722, x_2723, x_2724, x_2725, x_2726, x_2727, x_2728, x_2729, x_2730, x_2731, x_2732, x_2733, x_2734, x_2735, x_2736, x_2737, x_2738, x_2739, x_2740, x_2741, x_2742, x_2743, x_2744, x_2745, x_2746, x_2747, x_2748, x_2749, x_2750, x_2751, x_2752, x_2753, x_2754, x_2755, x_2756, x_2757, x_2758, x_2759, x_2760, x_2761, x_2762, x_2763, x_2764, x_2765, x_2766, x_2767, x_2768, x_2769, x_2770, x_2771, x_2772, x_2773, x_2774, x_2775, x_2776, x_2777, x_2778, x_2779, x_2780, x_2781, x_2782, x_2783, x_2784, x_2785, x_2786, x_2787, x_2788, x_2789, x_2790, x_2791, x_2792, x_2793, x_2794, x_2795, x_2796, x_2797, x_2798, x_2799, x_2800, x_2801, x_2802, x_2803, x_2804, x_2805, x_2806, x_2807, x_2808, x_2809, x_2810, x_2811, x_2812, x_2813, x_2814, x_2815, x_2816, x_2817, x_2818, x_2819, x_2820, x_2821, x_2822, x_2823, x_2824, x_2825, x_2826, x_2827, x_2828, x_2829, x_2830, x_2831, x_2832, x_2833, x_2834, x_2835, x_2836, x_2837, x_2838, x_2839, x_2840, x_2841, x_2842, x_2843, x_2844, x_2845, x_2846, x_2847, x_2848, x_2849, x_2850, x_2851, x_2852, x_2853, x_2854, x_2855, x_2856, x_2857, x_2858, x_2859, x_2860, x_2861, x_2862, x_2863, x_2864, x_2865, x_2866, x_2867, x_2868, x_2869, x_2870, x_2871, x_2872, x_2873, x_2874, x_2875, x_2876, x_2877, x_2878, x_2879, x_2880, x_2881, x_2882, x_2883, x_2884, x_2885, x_2886, x_2887, x_2888, x_2889, x_2890, x_2891, x_2892, x_2893, x_2894, x_2895, x_2896, x_2897, x_2898, x_2899, x_2900, x_2901, x_2902, x_2903, x_2904, x_2905, x_2906, x_2907, x_2908, x_2909, x_2910, x_2911, x_2912, x_2913, x_2914, x_2915, x_2916, x_2917, x_2918, x_2919, x_2920, x_2921, x_2922, x_2923, x_2924, x_2925, x_2926, x_2927, x_2928, x_2929, x_2930, x_2931, x_2932, x_2933, x_2934, x_2935, x_2936, x_2937, x_2938, x_2939, x_2940, x_2941, x_2942, x_2943, x_2944, x_2945, x_2946, x_2947, x_2948, x_2949, x_2950, x_2951, x_2952, x_2953, x_2954, x_2955, x_2956, x_2957, x_2958, x_2959, x_2960, x_2961, x_2962, x_2963, x_2964, x_2965, x_2966, x_2967, x_2968, x_2969, x_2970, x_2971, x_2972, x_2973, x_2974, x_2975, x_2976, x_2977, x_2978, x_2979, x_2980, x_2981, x_2982, x_2983, x_2984, x_2985, x_2986, x_2987, x_2988, x_2989, x_2990, x_2991, x_2992, x_2993, x_2994, x_2995, x_2996, x_2997, x_2998, x_2999, x_3000, x_3001, x_3002, x_3003, x_3004, x_3005, x_3006, x_3007, x_3008, x_3009, x_3010, x_3011, x_3012, x_3013, x_3014, x_3015, x_3016, x_3017, x_3018, x_3019, x_3020, x_3021, x_3022, x_3023, x_3024, x_3025, x_3026, x_3027, x_3028, x_3029, x_3030, x_3031, x_3032, x_3033, x_3034, x_3035, x_3036, x_3037, x_3038, x_3039, x_3040, x_3041, x_3042, x_3043, x_3044, x_3045, x_3046, x_3047, x_3048, x_3049, x_3050, x_3051, x_3052, x_3053, x_3054, x_3055, x_3056, x_3057, x_3058, x_3059, x_3060, x_3061, x_3062, x_3063, x_3064, x_3065, x_3066, x_3067, x_3068, x_3069, x_3070, x_3071, x_3072, x_3073, x_3074, x_3075, x_3076, x_3077, x_3078, x_3079, x_3080, x_3081, x_3082, x_3083, x_3084, x_3085, x_3086, x_3087, x_3088, x_3089, x_3090, x_3091, x_3092, x_3093, x_3094, x_3095, x_3096, x_3097, x_3098, x_3099, x_3100, x_3101, x_3102, x_3103, x_3104, x_3105, x_3106, x_3107, x_3108, x_3109, x_3110, x_3111, x_3112, x_3113, x_3114, x_3115, x_3116, x_3117, x_3118, x_3119, x_3120, x_3121, x_3122, x_3123, x_3124, x_3125, x_3126, x_3127, x_3128, x_3129, x_3130, x_3131, x_3132, x_3133, x_3134, x_3135, x_3136, x_3137, x_3138, x_3139, x_3140, x_3141, x_3142, x_3143, x_3144, x_3145, x_3146, x_3147, x_3148, x_3149, x_3150, x_3151, x_3152, x_3153, x_3154, x_3155, x_3156, x_3157, x_3158, x_3159, x_3160, x_3161, x_3162, x_3163, x_3164, x_3165, x_3166, x_3167, x_3168, x_3169, x_3170, x_3171, x_3172, x_3173, x_3174, x_3175, x_3176, x_3177, x_3178, x_3179, x_3180, x_3181, x_3182, x_3183, x_3184, x_3185, x_3186, x_3187, x_3188, x_3189, x_3190, x_3191, x_3192, x_3193, x_3194, x_3195, x_3196, x_3197, x_3198, x_3199, x_3200, x_3201, x_3202, x_3203, x_3204, x_3205, x_3206, x_3207, x_3208, x_3209, x_3210, x_3211, x_3212, x_3213, x_3214, x_3215, x_3216, x_3217, x_3218, x_3219, x_3220, x_3221, x_3222, x_3223, x_3224, x_3225, x_3226, x_3227, x_3228, x_3229, x_3230, x_3231, x_3232, x_3233, x_3234, x_3235, x_3236, x_3237, x_3238, x_3239, x_3240, x_3241, x_3242, x_3243, x_3244, x_3245, x_3246, x_3247, x_3248, x_3249, x_3250, x_3251, x_3252, x_3253, x_3254, x_3255, x_3256, x_3257, x_3258, x_3259, x_3260, x_3261, x_3262, x_3263, x_3264, x_3265, x_3266, x_3267, x_3268, x_3269, x_3270, x_3271, x_3272, x_3273, x_3274, x_3275, x_3276, x_3277, x_3278, x_3279, x_3280, x_3281, x_3282, x_3283, x_3284, x_3285, x_3286, x_3287, x_3288, x_3289, x_3290, x_3291, x_3292, x_3293, x_3294, x_3295, x_3296, x_3297, x_3298, x_3299, x_3300, x_3301, x_3302, x_3303, x_3304, x_3305, x_3306, x_3307, x_3308, x_3309, x_3310, x_3311, x_3312, x_3313, x_3314, x_3315, x_3316, x_3317, x_3318, x_3319, x_3320, x_3321, x_3322, x_3323, x_3324, x_3325, x_3326, x_3327, x_3328, x_3329, x_3330, x_3331, x_3332, x_3333, x_3334, x_3335, x_3336, x_3337, x_3338, x_3339, x_3340, x_3341, x_3342, x_3343, x_3344, x_3345, x_3346, x_3347, x_3348, x_3349, x_3350, x_3351, x_3352, x_3353, x_3354, x_3355, x_3356, x_3357, x_3358, x_3359, x_3360, x_3361, x_3362, x_3363, x_3364, x_3365, x_3366, x_3367, x_3368, x_3369, x_3370, x_3371, x_3372, x_3373, x_3374, x_3375, x_3376, x_3377, x_3378, x_3379, x_3380, x_3381, x_3382, x_3383, x_3384, x_3385, x_3386, x_3387, x_3388, x_3389, x_3390, x_3391, x_3392, x_3393, x_3394, x_3395, x_3396, x_3397, x_3398, x_3399, x_3400, x_3401, x_3402, x_3403, x_3404, x_3405, x_3406, x_3407, x_3408, x_3409, x_3410, x_3411, x_3412, x_3413, x_3414, x_3415, x_3416, x_3417, x_3418, x_3419, x_3420, x_3421, x_3422, x_3423, x_3424, x_3425, x_3426, x_3427, x_3428, x_3429, x_3430, x_3431, x_3432, x_3433, x_3434, x_3435, x_3436, x_3437, x_3438, x_3439, x_3440, x_3441, x_3442, x_3443, x_3444, x_3445, x_3446, x_3447, x_3448, x_3449, x_3450, x_3451, x_3452, x_3453, x_3454, x_3455, x_3456, x_3457, x_3458, x_3459, x_3460, x_3461, x_3462, x_3463, x_3464, x_3465, x_3466, x_3467, x_3468, x_3469, x_3470, x_3471, x_3472, x_3473, x_3474, x_3475, x_3476, x_3477, x_3478, x_3479, x_3480, x_3481, x_3482, x_3483, x_3484, x_3485, x_3486, x_3487, x_3488, x_3489, x_3490, x_3491, x_3492, x_3493, x_3494, x_3495, x_3496, x_3497, x_3498, x_3499, x_3500, x_3501, x_3502, x_3503, x_3504, x_3505, x_3506, x_3507, x_3508, x_3509, x_3510, x_3511, x_3512, x_3513, x_3514, x_3515, x_3516, x_3517, x_3518, x_3519, x_3520, x_3521, x_3522, x_3523, x_3524, x_3525, x_3526, x_3527, x_3528, x_3529, x_3530, x_3531, x_3532, x_3533, x_3534, x_3535, x_3536, x_3537, x_3538, x_3539, x_3540, x_3541, x_3542, x_3543, x_3544, x_3545, x_3546, x_3547, x_3548, x_3549, x_3550, x_3551, x_3552, x_3553, x_3554, x_3555, x_3556, x_3557, x_3558, x_3559, x_3560, x_3561, x_3562, x_3563, x_3564, x_3565, x_3566, x_3567, x_3568, x_3569, x_3570, x_3571, x_3572, x_3573, x_3574, x_3575, x_3576, x_3577, x_3578, x_3579, x_3580, x_3581, x_3582, x_3583, x_3584, x_3585, x_3586, x_3587, x_3588, x_3589, x_3590, x_3591, x_3592, x_3593, x_3594, x_3595, x_3596, x_3597, x_3598, x_3599, x_3600, x_3601, x_3602, x_3603, x_3604, x_3605, x_3606, x_3607, x_3608, x_3609, x_3610, x_3611, x_3612, x_3613, x_3614, x_3615, x_3616, x_3617, x_3618, x_3619, x_3620, x_3621, x_3622, x_3623, x_3624, x_3625, x_3626, x_3627, x_3628, x_3629, x_3630, x_3631, x_3632, x_3633, x_3634, x_3635, x_3636, x_3637, x_3638, x_3639, x_3640, x_3641, x_3642, x_3643, x_3644, x_3645, x_3646, x_3647, x_3648, x_3649, x_3650, x_3651, x_3652, x_3653, x_3654, x_3655, x_3656, x_3657, x_3658, x_3659, x_3660, x_3661, x_3662, x_3663, x_3664, x_3665, x_3666, x_3667, x_3668, x_3669, x_3670, x_3671, x_3672, x_3673, x_3674, x_3675, x_3676, x_3677, x_3678, x_3679, x_3680, x_3681, x_3682, x_3683, x_3684, x_3685, x_3686, x_3687, x_3688, x_3689, x_3690, x_3691, x_3692, x_3693, x_3694, x_3695, x_3696, x_3697, x_3698, x_3699, x_3700, x_3701, x_3702, x_3703, x_3704, x_3705, x_3706, x_3707, x_3708, x_3709, x_3710, x_3711, x_3712, x_3713, x_3714, x_3715, x_3716, x_3717, x_3718, x_3719, x_3720, x_3721, x_3722, x_3723, x_3724, x_3725, x_3726, x_3727, x_3728, x_3729, x_3730, x_3731, x_3732, x_3733, x_3734, x_3735, x_3736, x_3737, x_3738, x_3739, x_3740, x_3741, x_3742, x_3743, x_3744, x_3745, x_3746, x_3747, x_3748, x_3749, x_3750, x_3751, x_3752, x_3753, x_3754, x_3755, x_3756, x_3757, x_3758, x_3759, x_3760, x_3761, x_3762, x_3763, x_3764, x_3765, x_3766, x_3767, x_3768, x_3769, x_3770, x_3771, x_3772, x_3773, x_3774, x_3775, x_3776, x_3777, x_3778, x_3779, x_3780, x_3781, x_3782, x_3783, x_3784, x_3785, x_3786, x_3787, x_3788, x_3789, x_3790, x_3791, x_3792, x_3793, x_3794, x_3795, x_3796, x_3797, x_3798, x_3799, x_3800, x_3801, x_3802, x_3803, x_3804, x_3805, x_3806, x_3807, x_3808, x_3809, x_3810, x_3811, x_3812, x_3813, x_3814, x_3815, x_3816, x_3817, x_3818, x_3819, x_3820, x_3821, x_3822, x_3823, x_3824, x_3825, x_3826, x_3827, x_3828, x_3829, x_3830, x_3831, x_3832, x_3833, x_3834, x_3835, x_3836, x_3837, x_3838, x_3839, x_3840, x_3841, x_3842, x_3843, x_3844, x_3845, x_3846, x_3847, x_3848, x_3849, x_3850, x_3851, x_3852, x_3853, x_3854, x_3855, x_3856, x_3857, x_3858, x_3859, x_3860, x_3861, x_3862, x_3863, x_3864, x_3865, x_3866, x_3867, x_3868, x_3869, x_3870, x_3871, x_3872, x_3873, x_3874, x_3875, x_3876, x_3877, x_3878, x_3879, x_3880, x_3881, x_3882, x_3883, x_3884, x_3885, x_3886, x_3887, x_3888, x_3889, x_3890, x_3891, x_3892, x_3893, x_3894, x_3895, x_3896, x_3897, x_3898, x_3899, x_3900, x_3901, x_3902, x_3903, x_3904, x_3905, x_3906, x_3907, x_3908, x_3909, x_3910, x_3911, x_3912, x_3913, x_3914, x_3915, x_3916, x_3917, x_3918, x_3919, x_3920, x_3921, x_3922, x_3923, x_3924, x_3925, x_3926, x_3927, x_3928, x_3929, x_3930, x_3931, x_3932, x_3933, x_3934, x_3935, x_3936, x_3937, x_3938, x_3939, x_3940, x_3941, x_3942, x_3943, x_3944, x_3945, x_3946, x_3947, x_3948, x_3949, x_3950, x_3951, x_3952, x_3953, x_3954, x_3955, x_3956, x_3957, x_3958, x_3959, x_3960, x_3961, x_3962, x_3963, x_3964, x_3965, x_3966, x_3967, x_3968, x_3969, x_3970, x_3971, x_3972, x_3973, x_3974, x_3975, x_3976, x_3977, x_3978, x_3979, x_3980, x_3981, x_3982, x_3983, x_3984, x_3985, x_3986, x_3987, x_3988, x_3989, x_3990, x_3991, x_3992, x_3993, x_3994, x_3995, x_3996, x_3997, x_3998, x_3999, x_4000, x_4001, x_4002, x_4003, x_4004, x_4005, x_4006, x_4007, x_4008, x_4009, x_4010, x_4011, x_4012, x_4013, x_4014, x_4015, x_4016, x_4017, x_4018, x_4019, x_4020, x_4021, x_4022, x_4023, x_4024, x_4025, x_4026, x_4027, x_4028, x_4029, x_4030, x_4031, x_4032, x_4033, x_4034, x_4035, x_4036, x_4037, x_4038, x_4039, x_4040, x_4041, x_4042, x_4043, x_4044, x_4045, x_4046, x_4047, x_4048, x_4049, x_4050, x_4051, x_4052, x_4053, x_4054, x_4055, x_4056, x_4057, x_4058, x_4059, x_4060, x_4061, x_4062, x_4063, x_4064, x_4065, x_4066, x_4067, x_4068, x_4069, x_4070, x_4071, x_4072, x_4073, x_4074, x_4075, x_4076, x_4077, x_4078, x_4079, x_4080, x_4081, x_4082, x_4083, x_4084, x_4085, x_4086, x_4087, x_4088, x_4089, x_4090, x_4091, x_4092, x_4093, x_4094, x_4095, x_4096, x_4097, x_4098, x_4099, x_4100, x_4101, x_4102, x_4103, x_4104, x_4105, x_4106, x_4107, x_4108, x_4109, x_4110, x_4111, x_4112, x_4113, x_4114, x_4115, x_4116, x_4117, x_4118, x_4119, x_4120, x_4121, x_4122, x_4123, x_4124, x_4125, x_4126, x_4127, x_4128, x_4129, x_4130, x_4131, x_4132, x_4133, x_4134, x_4135, x_4136, x_4137, x_4138, x_4139, x_4140, x_4141, x_4142, x_4143, x_4144, x_4145, x_4146, x_4147, x_4148, x_4149, x_4150, x_4151, x_4152, x_4153, x_4154, x_4155, x_4156, x_4157, x_4158, x_4159, x_4160, x_4161, x_4162, x_4163, x_4164, x_4165, x_4166, x_4167, x_4168, x_4169, x_4170, x_4171, x_4172, x_4173, x_4174, x_4175, x_4176, x_4177, x_4178, x_4179, x_4180, x_4181, x_4182, x_4183, x_4184, x_4185, x_4186, x_4187, x_4188, x_4189, x_4190, x_4191, x_4192, x_4193, x_4194, x_4195, x_4196, x_4197, x_4198, x_4199, x_4200, x_4201, x_4202, x_4203, x_4204, x_4205, x_4206, x_4207, x_4208, x_4209, x_4210, x_4211, x_4212, x_4213, x_4214, x_4215, x_4216, x_4217, x_4218, x_4219, x_4220, x_4221, x_4222, x_4223, x_4224, x_4225, x_4226, x_4227, x_4228, x_4229, x_4230, x_4231, x_4232, x_4233, x_4234, x_4235, x_4236, x_4237, x_4238, x_4239, x_4240, x_4241, x_4242, x_4243, x_4244, x_4245, x_4246, x_4247, x_4248, x_4249, x_4250, x_4251, x_4252, x_4253, x_4254, x_4255, x_4256, x_4257, x_4258, x_4259, x_4260, x_4261, x_4262, x_4263, x_4264, x_4265, x_4266, x_4267, x_4268, x_4269, x_4270, x_4271, x_4272, x_4273, x_4274, x_4275, x_4276, x_4277, x_4278, x_4279, x_4280, x_4281, x_4282, x_4283, x_4284, x_4285, x_4286, x_4287, x_4288, x_4289, x_4290, x_4291, x_4292, x_4293, x_4294, x_4295, x_4296, x_4297, x_4298, x_4299, x_4300, x_4301, x_4302, x_4303, x_4304, x_4305, x_4306, x_4307, x_4308, x_4309, x_4310, x_4311, x_4312, x_4313, x_4314, x_4315, x_4316, x_4317, x_4318, x_4319, x_4320, x_4321, x_4322, x_4323, x_4324, x_4325, x_4326, x_4327, x_4328, x_4329, x_4330, x_4331, x_4332, x_4333, x_4334, x_4335, x_4336, x_4337, x_4338, x_4339, x_4340, x_4341, x_4342, x_4343, x_4344, x_4345, x_4346, x_4347, x_4348, x_4349, x_4350, x_4351, x_4352, x_4353, x_4354, x_4355, x_4356, x_4357, x_4358, x_4359, x_4360, x_4361, x_4362, x_4363, x_4364, x_4365, x_4366, x_4367, x_4368, x_4369, x_4370, x_4371, x_4372, x_4373, x_4374, x_4375, x_4376, x_4377, x_4378, x_4379, x_4380, x_4381, x_4382, x_4383, x_4384, x_4385, x_4386, x_4387, x_4388, x_4389, x_4390, x_4391, x_4392, x_4393, x_4394, x_4395, x_4396, x_4397, x_4398, x_4399, x_4400, x_4401, x_4402, x_4403, x_4404, x_4405, x_4406, x_4407, x_4408, x_4409, x_4410, x_4411, x_4412, x_4413, x_4414, x_4415, x_4416, x_4417, x_4418, x_4419, x_4420, x_4421, x_4422, x_4423, x_4424, x_4425, x_4426, x_4427, x_4428, x_4429, x_4430, x_4431, x_4432, x_4433, x_4434, x_4435, x_4436, x_4437, x_4438, x_4439, x_4440, x_4441, x_4442, x_4443, x_4444, x_4445, x_4446, x_4447, x_4448, x_4449, x_4450, x_4451, x_4452, x_4453, x_4454, x_4455, x_4456, x_4457, x_4458, x_4459, x_4460, x_4461, x_4462, x_4463, x_4464, x_4465, x_4466, x_4467, x_4468, x_4469, x_4470, x_4471, x_4472, x_4473, x_4474, x_4475, x_4476, x_4477, x_4478, x_4479, x_4480, x_4481, x_4482, x_4483, x_4484, x_4485, x_4486, x_4487, x_4488, x_4489, x_4490, x_4491, x_4492, x_4493, x_4494, x_4495, x_4496, x_4497, x_4498, x_4499, x_4500, x_4501, x_4502, x_4503, x_4504, x_4505, x_4506, x_4507, x_4508, x_4509, x_4510, x_4511, x_4512, x_4513, x_4514, x_4515, x_4516, x_4517, x_4518, x_4519, x_4520, x_4521, x_4522, x_4523, x_4524, x_4525, x_4526, x_4527, x_4528, x_4529, x_4530, x_4531, x_4532, x_4533, x_4534, x_4535, x_4536, x_4537, x_4538, x_4539, x_4540, x_4541, x_4542, x_4543, x_4544, x_4545, x_4546, x_4547, x_4548, x_4549, x_4550, x_4551, x_4552, x_4553, x_4554, x_4555, x_4556, x_4557, x_4558, x_4559, x_4560, x_4561, x_4562, x_4563, x_4564, x_4565, x_4566, x_4567, x_4568, x_4569, x_4570, x_4571, x_4572, x_4573, x_4574, x_4575, x_4576, x_4577, x_4578, x_4579, x_4580, x_4581, x_4582, x_4583, x_4584, x_4585, x_4586, x_4587, x_4588, x_4589, x_4590, x_4591, x_4592, x_4593, x_4594, x_4595, x_4596, x_4597, x_4598, x_4599, x_4600, x_4601, x_4602, x_4603, x_4604, x_4605, x_4606, x_4607, x_4608, x_4609, x_4610, x_4611, x_4612, x_4613, x_4614, x_4615, x_4616, x_4617, x_4618, x_4619, x_4620, x_4621, x_4622, x_4623, x_4624, x_4625, x_4626, x_4627, x_4628, x_4629, x_4630, x_4631, x_4632, x_4633, x_4634, x_4635, x_4636, x_4637, x_4638, x_4639, x_4640, x_4641, x_4642, x_4643, x_4644, x_4645, x_4646, x_4647, x_4648, x_4649, x_4650, x_4651, x_4652, x_4653, x_4654, x_4655, x_4656, x_4657, x_4658, x_4659, x_4660, x_4661, x_4662, x_4663, x_4664, x_4665, x_4666, x_4667, x_4668, x_4669, x_4670, x_4671, x_4672, x_4673, x_4674, x_4675, x_4676, x_4677, x_4678, x_4679, x_4680, x_4681, x_4682, x_4683, x_4684, x_4685, x_4686, x_4687, x_4688, x_4689, x_4690, x_4691, x_4692, x_4693, x_4694, x_4695, x_4696, x_4697, x_4698, x_4699, x_4700, x_4701, x_4702, x_4703, x_4704, x_4705, x_4706, x_4707, x_4708, x_4709, x_4710, x_4711, x_4712, x_4713, x_4714, x_4715, x_4716, x_4717, x_4718, x_4719, x_4720, x_4721, x_4722, x_4723, x_4724, x_4725, x_4726, x_4727, x_4728, x_4729, x_4730, x_4731, x_4732, x_4733, x_4734, x_4735, x_4736, x_4737, x_4738, x_4739, x_4740, x_4741, x_4742, x_4743, x_4744, x_4745, x_4746, x_4747, x_4748, x_4749, x_4750, x_4751, x_4752, x_4753, x_4754, x_4755, x_4756, x_4757, x_4758, x_4759, x_4760, x_4761, x_4762, x_4763, x_4764, x_4765, x_4766, x_4767, x_4768, x_4769, x_4770, x_4771, x_4772, x_4773, x_4774, x_4775, x_4776, x_4777, x_4778, x_4779, x_4780, x_4781, x_4782, x_4783, x_4784, x_4785, x_4786, x_4787, x_4788, x_4789, x_4790, x_4791, x_4792, x_4793, x_4794, x_4795, x_4796, x_4797, x_4798, x_4799, x_4800, x_4801, x_4802, x_4803, x_4804, x_4805, x_4806, x_4807, x_4808, x_4809, x_4810, x_4811, x_4812, x_4813, x_4814, x_4815, x_4816, x_4817, x_4818, x_4819, x_4820, x_4821, x_4822, x_4823, x_4824, x_4825, x_4826, x_4827, x_4828, x_4829, x_4830, x_4831, x_4832, x_4833, x_4834, x_4835, x_4836, x_4837, x_4838, x_4839, x_4840, x_4841, x_4842, x_4843, x_4844, x_4845, x_4846, x_4847, x_4848, x_4849, x_4850, x_4851, x_4852, x_4853, x_4854, x_4855, x_4856, x_4857, x_4858, x_4859, x_4860, x_4861, x_4862, x_4863, x_4864, x_4865, x_4866, x_4867, x_4868, x_4869, x_4870, x_4871, x_4872, x_4873, x_4874, x_4875, x_4876, x_4877, x_4878, x_4879, x_4880, x_4881, x_4882, x_4883, x_4884, x_4885, x_4886, x_4887, x_4888, x_4889, x_4890, x_4891, x_4892, x_4893, x_4894, x_4895, x_4896, x_4897, x_4898, x_4899, x_4900, x_4901, x_4902, x_4903, x_4904, x_4905, x_4906, x_4907, x_4908, x_4909, x_4910, x_4911, x_4912, x_4913, x_4914, x_4915, x_4916, x_4917, x_4918, x_4919, x_4920, x_4921, x_4922, x_4923, x_4924, x_4925, x_4926, x_4927, x_4928, x_4929, x_4930, x_4931, x_4932, x_4933, x_4934, x_4935, x_4936, x_4937, x_4938, x_4939, x_4940, x_4941, x_4942, x_4943, x_4944, x_4945, x_4946, x_4947, x_4948, x_4949, x_4950, x_4951, x_4952, x_4953, x_4954, x_4955, x_4956, x_4957, x_4958, x_4959, x_4960, x_4961, x_4962, x_4963, x_4964, x_4965, x_4966, x_4967, x_4968, x_4969, x_4970, x_4971, x_4972, x_4973, x_4974, x_4975, x_4976, x_4977, x_4978, x_4979, x_4980, x_4981, x_4982, x_4983, x_4984, x_4985, x_4986, x_4987, x_4988, x_4989, x_4990, x_4991, x_4992, x_4993, x_4994, x_4995, x_4996, x_4997, x_4998, x_4999, x_5000, x_5001, x_5002, x_5003, x_5004, x_5005, x_5006, x_5007, x_5008, x_5009, x_5010, x_5011, x_5012, x_5013, x_5014, x_5015, x_5016, x_5017, x_5018, x_5019, x_5020, x_5021, x_5022, x_5023, x_5024, x_5025, x_5026, x_5027, x_5028, x_5029, x_5030, x_5031, x_5032, x_5033, x_5034, x_5035, x_5036, x_5037, x_5038, x_5039, x_5040, x_5041, x_5042, x_5043, x_5044, x_5045, x_5046, x_5047, x_5048, x_5049, x_5050, x_5051, x_5052, x_5053, x_5054, x_5055, x_5056, x_5057, x_5058, x_5059, x_5060, x_5061, x_5062, x_5063, x_5064, x_5065, x_5066, x_5067, x_5068, x_5069, x_5070, x_5071, x_5072, x_5073, x_5074, x_5075, x_5076, x_5077, x_5078, x_5079, x_5080, x_5081, x_5082, x_5083, x_5084, x_5085, x_5086, x_5087, x_5088, x_5089, x_5090, x_5091, x_5092, x_5093, x_5094, x_5095, x_5096, x_5097, x_5098, x_5099, x_5100, x_5101, x_5102, x_5103, x_5104, x_5105, x_5106, x_5107, x_5108, x_5109, x_5110, x_5111, x_5112, x_5113, x_5114, x_5115, x_5116, x_5117, x_5118, x_5119, x_5120, x_5121, x_5122, x_5123, x_5124, x_5125, x_5126, x_5127, x_5128, x_5129, x_5130, x_5131, x_5132, x_5133, x_5134, x_5135, x_5136, x_5137, x_5138, x_5139, x_5140, x_5141, x_5142, x_5143, x_5144, x_5145, x_5146, x_5147, x_5148, x_5149, x_5150, x_5151, x_5152, x_5153, x_5154, x_5155, x_5156, x_5157, x_5158, x_5159, x_5160, x_5161, x_5162, x_5163, x_5164, x_5165, x_5166, x_5167, x_5168, x_5169, x_5170, x_5171, x_5172, x_5173, x_5174, x_5175, x_5176, x_5177, x_5178, x_5179, x_5180, x_5181, x_5182, x_5183, x_5184, x_5185, x_5186, x_5187, x_5188, x_5189, x_5190, x_5191, x_5192, x_5193, x_5194, x_5195, x_5196, x_5197, x_5198, x_5199, x_5200, x_5201, x_5202, x_5203, x_5204, x_5205, x_5206, x_5207, x_5208, x_5209, x_5210, x_5211, x_5212, x_5213, x_5214, x_5215, x_5216, x_5217, x_5218, x_5219, x_5220, x_5221, x_5222, x_5223, x_5224, x_5225, x_5226, x_5227, x_5228, x_5229, x_5230, x_5231, x_5232, x_5233, x_5234, x_5235, x_5236, x_5237, x_5238, x_5239, x_5240, x_5241, x_5242, x_5243, x_5244, x_5245, x_5246, x_5247, x_5248, x_5249, x_5250, x_5251, x_5252, x_5253, x_5254, x_5255, x_5256, x_5257, x_5258, x_5259, x_5260, x_5261, x_5262, x_5263, x_5264, x_5265, x_5266, x_5267, x_5268, x_5269, x_5270, x_5271, x_5272, x_5273, x_5274, x_5275, x_5276, x_5277, x_5278, x_5279, x_5280, x_5281, x_5282, x_5283, x_5284, x_5285, x_5286, x_5287, x_5288, x_5289, x_5290, x_5291, x_5292, x_5293, x_5294, x_5295, x_5296, x_5297, x_5298, x_5299, x_5300, x_5301, x_5302, x_5303, x_5304, x_5305, x_5306, x_5307, x_5308, x_5309, x_5310, x_5311, x_5312, x_5313, x_5314, x_5315, x_5316, x_5317, x_5318, x_5319, x_5320, x_5321, x_5322, x_5323, x_5324, x_5325, x_5326, x_5327, x_5328, x_5329, x_5330, x_5331, x_5332, x_5333, x_5334, x_5335, x_5336, x_5337, x_5338, x_5339, x_5340, x_5341, x_5342, x_5343, x_5344, x_5345, x_5346, x_5347, x_5348, x_5349, x_5350, x_5351, x_5352, x_5353, x_5354, x_5355, x_5356, x_5357, x_5358, x_5359, x_5360, x_5361, x_5362, x_5363, x_5364, x_5365, x_5366, x_5367, x_5368, x_5369, x_5370, x_5371, x_5372, x_5373, x_5374, x_5375, x_5376, x_5377, x_5378, x_5379, x_5380, x_5381, x_5382, x_5383, x_5384, x_5385, x_5386, x_5387, x_5388, x_5389, x_5390, x_5391, x_5392, x_5393, x_5394, x_5395, x_5396, x_5397, x_5398, x_5399, x_5400, x_5401, x_5402, x_5403, x_5404, x_5405, x_5406, x_5407, x_5408, x_5409, x_5410, x_5411, x_5412, x_5413, x_5414, x_5415, x_5416, x_5417, x_5418, x_5419, x_5420, x_5421, x_5422, x_5423, x_5424, x_5425, x_5426, x_5427, x_5428, x_5429, x_5430, x_5431, x_5432, x_5433, x_5434, x_5435, x_5436, x_5437, x_5438, x_5439, x_5440, x_5441, x_5442, x_5443, x_5444, x_5445, x_5446, x_5447, x_5448, x_5449, x_5450, x_5451, x_5452, x_5453, x_5454, x_5455, x_5456, x_5457, x_5458, x_5459, x_5460, x_5461, x_5462, x_5463, x_5464, x_5465, x_5466, x_5467, x_5468, x_5469, x_5470, x_5471, x_5472, x_5473, x_5474, x_5475, x_5476, x_5477, x_5478, x_5479, x_5480, x_5481, x_5482, x_5483, x_5484, x_5485, x_5486, x_5487, x_5488, x_5489, x_5490, x_5491, x_5492, x_5493, x_5494, x_5495, x_5496, x_5497, x_5498, x_5499, x_5500, x_5501, x_5502, x_5503, x_5504, x_5505, x_5506, x_5507, x_5508, x_5509, x_5510, x_5511, x_5512, x_5513, x_5514, x_5515, x_5516, x_5517, x_5518, x_5519, x_5520, x_5521, x_5522, x_5523, x_5524, x_5525, x_5526, x_5527, x_5528, x_5529, x_5530, x_5531, x_5532, x_5533, x_5534, x_5535, x_5536, x_5537, x_5538, x_5539, x_5540, x_5541, x_5542, x_5543, x_5544, x_5545, x_5546, x_5547, x_5548, x_5549, x_5550, x_5551, x_5552, x_5553, x_5554, x_5555, x_5556, x_5557, x_5558, x_5559, x_5560, x_5561, x_5562, x_5563, x_5564, x_5565, x_5566, x_5567, x_5568, x_5569, x_5570, x_5571, x_5572, x_5573, x_5574, x_5575, x_5576, x_5577, x_5578, x_5579, x_5580, x_5581, x_5582, x_5583, x_5584, x_5585, x_5586, x_5587, x_5588, x_5589, x_5590, x_5591, x_5592, x_5593, x_5594, x_5595, x_5596, x_5597, x_5598, x_5599, x_5600, x_5601, x_5602, x_5603, x_5604, x_5605, x_5606, x_5607, x_5608, x_5609, x_5610, x_5611, x_5612, x_5613, x_5614, x_5615, x_5616, x_5617, x_5618, x_5619, x_5620, x_5621, x_5622, x_5623, x_5624, x_5625, x_5626, x_5627, x_5628, x_5629, x_5630, x_5631, x_5632, x_5633, x_5634, x_5635, x_5636, x_5637, x_5638, x_5639, x_5640, x_5641, x_5642, x_5643, x_5644, x_5645, x_5646, x_5647, x_5648, x_5649, x_5650, x_5651, x_5652, x_5653, x_5654, x_5655, x_5656, x_5657, x_5658, x_5659, x_5660, x_5661, x_5662, x_5663, x_5664, x_5665, x_5666, x_5667, x_5668, x_5669, x_5670, x_5671, x_5672, x_5673, x_5674, x_5675, x_5676, x_5677, x_5678, x_5679, x_5680, x_5681, x_5682, x_5683, x_5684, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input x_33;
input x_34;
input x_35;
input x_36;
input x_37;
input x_38;
input x_39;
input x_40;
input x_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
input x_181;
input x_182;
input x_183;
input x_184;
input x_185;
input x_186;
input x_187;
input x_188;
input x_189;
input x_190;
input x_191;
input x_192;
input x_193;
input x_194;
input x_195;
input x_196;
input x_197;
input x_198;
input x_199;
input x_200;
input x_201;
input x_202;
input x_203;
input x_204;
input x_205;
input x_206;
input x_207;
input x_208;
input x_209;
input x_210;
input x_211;
input x_212;
input x_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
input x_460;
input x_461;
input x_462;
input x_463;
input x_464;
input x_465;
input x_466;
input x_467;
input x_468;
input x_469;
input x_470;
input x_471;
input x_472;
input x_473;
input x_474;
input x_475;
input x_476;
input x_477;
input x_478;
input x_479;
input x_480;
input x_481;
input x_482;
input x_483;
input x_484;
input x_485;
input x_486;
input x_487;
input x_488;
input x_489;
input x_490;
input x_491;
input x_492;
input x_493;
input x_494;
input x_495;
input x_496;
input x_497;
input x_498;
input x_499;
input x_500;
input x_501;
input x_502;
input x_503;
input x_504;
input x_505;
input x_506;
input x_507;
input x_508;
input x_509;
input x_510;
input x_511;
input x_512;
input x_513;
input x_514;
input x_515;
input x_516;
input x_517;
input x_518;
input x_519;
input x_520;
input x_521;
input x_522;
input x_523;
input x_524;
input x_525;
input x_526;
input x_527;
input x_528;
input x_529;
input x_530;
input x_531;
input x_532;
input x_533;
input x_534;
input x_535;
input x_536;
input x_537;
input x_538;
input x_539;
input x_540;
input x_541;
input x_542;
input x_543;
input x_544;
input x_545;
input x_546;
input x_547;
input x_548;
input x_549;
input x_550;
input x_551;
input x_552;
input x_553;
input x_554;
input x_555;
input x_556;
input x_557;
input x_558;
input x_559;
input x_560;
input x_561;
input x_562;
input x_563;
input x_564;
input x_565;
input x_566;
input x_567;
input x_568;
input x_569;
input x_570;
input x_571;
input x_572;
input x_573;
input x_574;
input x_575;
input x_576;
input x_577;
input x_578;
input x_579;
input x_580;
input x_581;
input x_582;
input x_583;
input x_584;
input x_585;
input x_586;
input x_587;
input x_588;
input x_589;
input x_590;
input x_591;
input x_592;
input x_593;
input x_594;
input x_595;
input x_596;
input x_597;
input x_598;
input x_599;
input x_600;
input x_601;
input x_602;
input x_603;
input x_604;
input x_605;
input x_606;
input x_607;
input x_608;
input x_609;
input x_610;
input x_611;
input x_612;
input x_613;
input x_614;
input x_615;
input x_616;
input x_617;
input x_618;
input x_619;
input x_620;
input x_621;
input x_622;
input x_623;
input x_624;
input x_625;
input x_626;
input x_627;
input x_628;
input x_629;
input x_630;
input x_631;
input x_632;
input x_633;
input x_634;
input x_635;
input x_636;
input x_637;
input x_638;
input x_639;
input x_640;
input x_641;
input x_642;
input x_643;
input x_644;
input x_645;
input x_646;
input x_647;
input x_648;
input x_649;
input x_650;
input x_651;
input x_652;
input x_653;
input x_654;
input x_655;
input x_656;
input x_657;
input x_658;
input x_659;
input x_660;
input x_661;
input x_662;
input x_663;
input x_664;
input x_665;
input x_666;
input x_667;
input x_668;
input x_669;
input x_670;
input x_671;
input x_672;
input x_673;
input x_674;
input x_675;
input x_676;
input x_677;
input x_678;
input x_679;
input x_680;
input x_681;
input x_682;
input x_683;
input x_684;
input x_685;
input x_686;
input x_687;
input x_688;
input x_689;
input x_690;
input x_691;
input x_692;
input x_693;
input x_694;
input x_695;
input x_696;
input x_697;
input x_698;
input x_699;
input x_700;
input x_701;
input x_702;
input x_703;
input x_704;
input x_705;
input x_706;
input x_707;
input x_708;
input x_709;
input x_710;
input x_711;
input x_712;
input x_713;
input x_714;
input x_715;
input x_716;
input x_717;
input x_718;
input x_719;
input x_720;
input x_721;
input x_722;
input x_723;
input x_724;
input x_725;
input x_726;
input x_727;
input x_728;
input x_729;
input x_730;
input x_731;
input x_732;
input x_733;
input x_734;
input x_735;
input x_736;
input x_737;
input x_738;
input x_739;
input x_740;
input x_741;
input x_742;
input x_743;
input x_744;
input x_745;
input x_746;
input x_747;
input x_748;
input x_749;
input x_750;
input x_751;
input x_752;
input x_753;
input x_754;
input x_755;
input x_756;
input x_757;
input x_758;
input x_759;
input x_760;
input x_761;
input x_762;
input x_763;
input x_764;
input x_765;
input x_766;
input x_767;
input x_768;
input x_769;
input x_770;
input x_771;
input x_772;
input x_773;
input x_774;
input x_775;
input x_776;
input x_777;
input x_778;
input x_779;
input x_780;
input x_781;
input x_782;
input x_783;
input x_784;
input x_785;
input x_786;
input x_787;
input x_788;
input x_789;
input x_790;
input x_791;
input x_792;
input x_793;
input x_794;
input x_795;
input x_796;
input x_797;
input x_798;
input x_799;
input x_800;
input x_801;
input x_802;
input x_803;
input x_804;
input x_805;
input x_806;
input x_807;
input x_808;
input x_809;
input x_810;
input x_811;
input x_812;
input x_813;
input x_814;
input x_815;
input x_816;
input x_817;
input x_818;
input x_819;
input x_820;
input x_821;
input x_822;
input x_823;
input x_824;
input x_825;
input x_826;
input x_827;
input x_828;
input x_829;
input x_830;
input x_831;
input x_832;
input x_833;
input x_834;
input x_835;
input x_836;
input x_837;
input x_838;
input x_839;
input x_840;
input x_841;
input x_842;
input x_843;
input x_844;
input x_845;
input x_846;
input x_847;
input x_848;
input x_849;
input x_850;
input x_851;
input x_852;
input x_853;
input x_854;
input x_855;
input x_856;
input x_857;
input x_858;
input x_859;
input x_860;
input x_861;
input x_862;
input x_863;
input x_864;
input x_865;
input x_866;
input x_867;
input x_868;
input x_869;
input x_870;
input x_871;
input x_872;
input x_873;
input x_874;
input x_875;
input x_876;
input x_877;
input x_878;
input x_879;
input x_880;
input x_881;
input x_882;
input x_883;
input x_884;
input x_885;
input x_886;
input x_887;
input x_888;
input x_889;
input x_890;
input x_891;
input x_892;
input x_893;
input x_894;
input x_895;
input x_896;
input x_897;
input x_898;
input x_899;
input x_900;
input x_901;
input x_902;
input x_903;
input x_904;
input x_905;
input x_906;
input x_907;
input x_908;
input x_909;
input x_910;
input x_911;
input x_912;
input x_913;
input x_914;
input x_915;
input x_916;
input x_917;
input x_918;
input x_919;
input x_920;
input x_921;
input x_922;
input x_923;
input x_924;
input x_925;
input x_926;
input x_927;
input x_928;
input x_929;
input x_930;
input x_931;
input x_932;
input x_933;
input x_934;
input x_935;
input x_936;
input x_937;
input x_938;
input x_939;
input x_940;
input x_941;
input x_942;
input x_943;
input x_944;
input x_945;
input x_946;
input x_947;
input x_948;
input x_949;
input x_950;
input x_951;
input x_952;
input x_953;
input x_954;
input x_955;
input x_956;
input x_957;
input x_958;
input x_959;
input x_960;
input x_961;
input x_962;
input x_963;
input x_964;
input x_965;
input x_966;
input x_967;
input x_968;
input x_969;
input x_970;
input x_971;
input x_972;
input x_973;
input x_974;
input x_975;
input x_976;
input x_977;
input x_978;
input x_979;
input x_980;
input x_981;
input x_982;
input x_983;
input x_984;
input x_985;
input x_986;
input x_987;
input x_988;
input x_989;
input x_990;
input x_991;
input x_992;
input x_993;
input x_994;
input x_995;
input x_996;
input x_997;
input x_998;
input x_999;
input x_1000;
input x_1001;
input x_1002;
input x_1003;
input x_1004;
input x_1005;
input x_1006;
input x_1007;
input x_1008;
input x_1009;
input x_1010;
input x_1011;
input x_1012;
input x_1013;
input x_1014;
input x_1015;
input x_1016;
input x_1017;
input x_1018;
input x_1019;
input x_1020;
input x_1021;
input x_1022;
input x_1023;
input x_1024;
input x_1025;
input x_1026;
input x_1027;
input x_1028;
input x_1029;
input x_1030;
input x_1031;
input x_1032;
input x_1033;
input x_1034;
input x_1035;
input x_1036;
input x_1037;
input x_1038;
input x_1039;
input x_1040;
input x_1041;
input x_1042;
input x_1043;
input x_1044;
input x_1045;
input x_1046;
input x_1047;
input x_1048;
input x_1049;
input x_1050;
input x_1051;
input x_1052;
input x_1053;
input x_1054;
input x_1055;
input x_1056;
input x_1057;
input x_1058;
input x_1059;
input x_1060;
input x_1061;
input x_1062;
input x_1063;
input x_1064;
input x_1065;
input x_1066;
input x_1067;
input x_1068;
input x_1069;
input x_1070;
input x_1071;
input x_1072;
input x_1073;
input x_1074;
input x_1075;
input x_1076;
input x_1077;
input x_1078;
input x_1079;
input x_1080;
input x_1081;
input x_1082;
input x_1083;
input x_1084;
input x_1085;
input x_1086;
input x_1087;
input x_1088;
input x_1089;
input x_1090;
input x_1091;
input x_1092;
input x_1093;
input x_1094;
input x_1095;
input x_1096;
input x_1097;
input x_1098;
input x_1099;
input x_1100;
input x_1101;
input x_1102;
input x_1103;
input x_1104;
input x_1105;
input x_1106;
input x_1107;
input x_1108;
input x_1109;
input x_1110;
input x_1111;
input x_1112;
input x_1113;
input x_1114;
input x_1115;
input x_1116;
input x_1117;
input x_1118;
input x_1119;
input x_1120;
input x_1121;
input x_1122;
input x_1123;
input x_1124;
input x_1125;
input x_1126;
input x_1127;
input x_1128;
input x_1129;
input x_1130;
input x_1131;
input x_1132;
input x_1133;
input x_1134;
input x_1135;
input x_1136;
input x_1137;
input x_1138;
input x_1139;
input x_1140;
input x_1141;
input x_1142;
input x_1143;
input x_1144;
input x_1145;
input x_1146;
input x_1147;
input x_1148;
input x_1149;
input x_1150;
input x_1151;
input x_1152;
input x_1153;
input x_1154;
input x_1155;
input x_1156;
input x_1157;
input x_1158;
input x_1159;
input x_1160;
input x_1161;
input x_1162;
input x_1163;
input x_1164;
input x_1165;
input x_1166;
input x_1167;
input x_1168;
input x_1169;
input x_1170;
input x_1171;
input x_1172;
input x_1173;
input x_1174;
input x_1175;
input x_1176;
input x_1177;
input x_1178;
input x_1179;
input x_1180;
input x_1181;
input x_1182;
input x_1183;
input x_1184;
input x_1185;
input x_1186;
input x_1187;
input x_1188;
input x_1189;
input x_1190;
input x_1191;
input x_1192;
input x_1193;
input x_1194;
input x_1195;
input x_1196;
input x_1197;
input x_1198;
input x_1199;
input x_1200;
input x_1201;
input x_1202;
input x_1203;
input x_1204;
input x_1205;
input x_1206;
input x_1207;
input x_1208;
input x_1209;
input x_1210;
input x_1211;
input x_1212;
input x_1213;
input x_1214;
input x_1215;
input x_1216;
input x_1217;
input x_1218;
input x_1219;
input x_1220;
input x_1221;
input x_1222;
input x_1223;
input x_1224;
input x_1225;
input x_1226;
input x_1227;
input x_1228;
input x_1229;
input x_1230;
input x_1231;
input x_1232;
input x_1233;
input x_1234;
input x_1235;
input x_1236;
input x_1237;
input x_1238;
input x_1239;
input x_1240;
input x_1241;
input x_1242;
input x_1243;
input x_1244;
input x_1245;
input x_1246;
input x_1247;
input x_1248;
input x_1249;
input x_1250;
input x_1251;
input x_1252;
input x_1253;
input x_1254;
input x_1255;
input x_1256;
input x_1257;
input x_1258;
input x_1259;
input x_1260;
input x_1261;
input x_1262;
input x_1263;
input x_1264;
input x_1265;
input x_1266;
input x_1267;
input x_1268;
input x_1269;
input x_1270;
input x_1271;
input x_1272;
input x_1273;
input x_1274;
input x_1275;
input x_1276;
input x_1277;
input x_1278;
input x_1279;
input x_1280;
input x_1281;
input x_1282;
input x_1283;
input x_1284;
input x_1285;
input x_1286;
input x_1287;
input x_1288;
input x_1289;
input x_1290;
input x_1291;
input x_1292;
input x_1293;
input x_1294;
input x_1295;
input x_1296;
input x_1297;
input x_1298;
input x_1299;
input x_1300;
input x_1301;
input x_1302;
input x_1303;
input x_1304;
input x_1305;
input x_1306;
input x_1307;
input x_1308;
input x_1309;
input x_1310;
input x_1311;
input x_1312;
input x_1313;
input x_1314;
input x_1315;
input x_1316;
input x_1317;
input x_1318;
input x_1319;
input x_1320;
input x_1321;
input x_1322;
input x_1323;
input x_1324;
input x_1325;
input x_1326;
input x_1327;
input x_1328;
input x_1329;
input x_1330;
input x_1331;
input x_1332;
input x_1333;
input x_1334;
input x_1335;
input x_1336;
input x_1337;
input x_1338;
input x_1339;
input x_1340;
input x_1341;
input x_1342;
input x_1343;
input x_1344;
input x_1345;
input x_1346;
input x_1347;
input x_1348;
input x_1349;
input x_1350;
input x_1351;
input x_1352;
input x_1353;
input x_1354;
input x_1355;
input x_1356;
input x_1357;
input x_1358;
input x_1359;
input x_1360;
input x_1361;
input x_1362;
input x_1363;
input x_1364;
input x_1365;
input x_1366;
input x_1367;
input x_1368;
input x_1369;
input x_1370;
input x_1371;
input x_1372;
input x_1373;
input x_1374;
input x_1375;
input x_1376;
input x_1377;
input x_1378;
input x_1379;
input x_1380;
input x_1381;
input x_1382;
input x_1383;
input x_1384;
input x_1385;
input x_1386;
input x_1387;
input x_1388;
input x_1389;
input x_1390;
input x_1391;
input x_1392;
input x_1393;
input x_1394;
input x_1395;
input x_1396;
input x_1397;
input x_1398;
input x_1399;
input x_1400;
input x_1401;
input x_1402;
input x_1403;
input x_1404;
input x_1405;
input x_1406;
input x_1407;
input x_1408;
input x_1409;
input x_1410;
input x_1411;
input x_1412;
input x_1413;
input x_1414;
input x_1415;
input x_1416;
input x_1417;
input x_1418;
input x_1419;
input x_1420;
input x_1421;
input x_1422;
input x_1423;
input x_1424;
input x_1425;
input x_1426;
input x_1427;
input x_1428;
input x_1429;
input x_1430;
input x_1431;
input x_1432;
input x_1433;
input x_1434;
input x_1435;
input x_1436;
input x_1437;
input x_1438;
input x_1439;
input x_1440;
input x_1441;
input x_1442;
input x_1443;
input x_1444;
input x_1445;
input x_1446;
input x_1447;
input x_1448;
input x_1449;
input x_1450;
input x_1451;
input x_1452;
input x_1453;
input x_1454;
input x_1455;
input x_1456;
input x_1457;
input x_1458;
input x_1459;
input x_1460;
input x_1461;
input x_1462;
input x_1463;
input x_1464;
input x_1465;
input x_1466;
input x_1467;
input x_1468;
input x_1469;
input x_1470;
input x_1471;
input x_1472;
input x_1473;
input x_1474;
input x_1475;
input x_1476;
input x_1477;
input x_1478;
input x_1479;
input x_1480;
input x_1481;
input x_1482;
input x_1483;
input x_1484;
input x_1485;
input x_1486;
input x_1487;
input x_1488;
input x_1489;
input x_1490;
input x_1491;
input x_1492;
input x_1493;
input x_1494;
input x_1495;
input x_1496;
input x_1497;
input x_1498;
input x_1499;
input x_1500;
input x_1501;
input x_1502;
input x_1503;
input x_1504;
input x_1505;
input x_1506;
input x_1507;
input x_1508;
input x_1509;
input x_1510;
input x_1511;
input x_1512;
input x_1513;
input x_1514;
input x_1515;
input x_1516;
input x_1517;
input x_1518;
input x_1519;
input x_1520;
input x_1521;
input x_1522;
input x_1523;
input x_1524;
input x_1525;
input x_1526;
input x_1527;
input x_1528;
input x_1529;
input x_1530;
input x_1531;
input x_1532;
input x_1533;
input x_1534;
input x_1535;
input x_1536;
input x_1537;
input x_1538;
input x_1539;
input x_1540;
input x_1541;
input x_1542;
input x_1543;
input x_1544;
input x_1545;
input x_1546;
input x_1547;
input x_1548;
input x_1549;
input x_1550;
input x_1551;
input x_1552;
input x_1553;
input x_1554;
input x_1555;
input x_1556;
input x_1557;
input x_1558;
input x_1559;
input x_1560;
input x_1561;
input x_1562;
input x_1563;
input x_1564;
input x_1565;
input x_1566;
input x_1567;
input x_1568;
input x_1569;
input x_1570;
input x_1571;
input x_1572;
input x_1573;
input x_1574;
input x_1575;
input x_1576;
input x_1577;
input x_1578;
input x_1579;
input x_1580;
input x_1581;
input x_1582;
input x_1583;
input x_1584;
input x_1585;
input x_1586;
input x_1587;
input x_1588;
input x_1589;
input x_1590;
input x_1591;
input x_1592;
input x_1593;
input x_1594;
input x_1595;
input x_1596;
input x_1597;
input x_1598;
input x_1599;
input x_1600;
input x_1601;
input x_1602;
input x_1603;
input x_1604;
input x_1605;
input x_1606;
input x_1607;
input x_1608;
input x_1609;
input x_1610;
input x_1611;
input x_1612;
input x_1613;
input x_1614;
input x_1615;
input x_1616;
input x_1617;
input x_1618;
input x_1619;
input x_1620;
input x_1621;
input x_1622;
input x_1623;
input x_1624;
input x_1625;
input x_1626;
input x_1627;
input x_1628;
input x_1629;
input x_1630;
input x_1631;
input x_1632;
input x_1633;
input x_1634;
input x_1635;
input x_1636;
input x_1637;
input x_1638;
input x_1639;
input x_1640;
input x_1641;
input x_1642;
input x_1643;
input x_1644;
input x_1645;
input x_1646;
input x_1647;
input x_1648;
input x_1649;
input x_1650;
input x_1651;
input x_1652;
input x_1653;
input x_1654;
input x_1655;
input x_1656;
input x_1657;
input x_1658;
input x_1659;
input x_1660;
input x_1661;
input x_1662;
input x_1663;
input x_1664;
input x_1665;
input x_1666;
input x_1667;
input x_1668;
input x_1669;
input x_1670;
input x_1671;
input x_1672;
input x_1673;
input x_1674;
input x_1675;
input x_1676;
input x_1677;
input x_1678;
input x_1679;
input x_1680;
input x_1681;
input x_1682;
input x_1683;
input x_1684;
input x_1685;
input x_1686;
input x_1687;
input x_1688;
input x_1689;
input x_1690;
input x_1691;
input x_1692;
input x_1693;
input x_1694;
input x_1695;
input x_1696;
input x_1697;
input x_1698;
input x_1699;
input x_1700;
input x_1701;
input x_1702;
input x_1703;
input x_1704;
input x_1705;
input x_1706;
input x_1707;
input x_1708;
input x_1709;
input x_1710;
input x_1711;
input x_1712;
input x_1713;
input x_1714;
input x_1715;
input x_1716;
input x_1717;
input x_1718;
input x_1719;
input x_1720;
input x_1721;
input x_1722;
input x_1723;
input x_1724;
input x_1725;
input x_1726;
input x_1727;
input x_1728;
input x_1729;
input x_1730;
input x_1731;
input x_1732;
input x_1733;
input x_1734;
input x_1735;
input x_1736;
input x_1737;
input x_1738;
input x_1739;
input x_1740;
input x_1741;
input x_1742;
input x_1743;
input x_1744;
input x_1745;
input x_1746;
input x_1747;
input x_1748;
input x_1749;
input x_1750;
input x_1751;
input x_1752;
input x_1753;
input x_1754;
input x_1755;
input x_1756;
input x_1757;
input x_1758;
input x_1759;
input x_1760;
input x_1761;
input x_1762;
input x_1763;
input x_1764;
input x_1765;
input x_1766;
input x_1767;
input x_1768;
input x_1769;
input x_1770;
input x_1771;
input x_1772;
input x_1773;
input x_1774;
input x_1775;
input x_1776;
input x_1777;
input x_1778;
input x_1779;
input x_1780;
input x_1781;
input x_1782;
input x_1783;
input x_1784;
input x_1785;
input x_1786;
input x_1787;
input x_1788;
input x_1789;
input x_1790;
input x_1791;
input x_1792;
input x_1793;
input x_1794;
input x_1795;
input x_1796;
input x_1797;
input x_1798;
input x_1799;
input x_1800;
input x_1801;
input x_1802;
input x_1803;
input x_1804;
input x_1805;
input x_1806;
input x_1807;
input x_1808;
input x_1809;
input x_1810;
input x_1811;
input x_1812;
input x_1813;
input x_1814;
input x_1815;
input x_1816;
input x_1817;
input x_1818;
input x_1819;
input x_1820;
input x_1821;
input x_1822;
input x_1823;
input x_1824;
input x_1825;
input x_1826;
input x_1827;
input x_1828;
input x_1829;
input x_1830;
input x_1831;
input x_1832;
input x_1833;
input x_1834;
input x_1835;
input x_1836;
input x_1837;
input x_1838;
input x_1839;
input x_1840;
input x_1841;
input x_1842;
input x_1843;
input x_1844;
input x_1845;
input x_1846;
input x_1847;
input x_1848;
input x_1849;
input x_1850;
input x_1851;
input x_1852;
input x_1853;
input x_1854;
input x_1855;
input x_1856;
input x_1857;
input x_1858;
input x_1859;
input x_1860;
input x_1861;
input x_1862;
input x_1863;
input x_1864;
input x_1865;
input x_1866;
input x_1867;
input x_1868;
input x_1869;
input x_1870;
input x_1871;
input x_1872;
input x_1873;
input x_1874;
input x_1875;
input x_1876;
input x_1877;
input x_1878;
input x_1879;
input x_1880;
input x_1881;
input x_1882;
input x_1883;
input x_1884;
input x_1885;
input x_1886;
input x_1887;
input x_1888;
input x_1889;
input x_1890;
input x_1891;
input x_1892;
input x_1893;
input x_1894;
input x_1895;
input x_1896;
input x_1897;
input x_1898;
input x_1899;
input x_1900;
input x_1901;
input x_1902;
input x_1903;
input x_1904;
input x_1905;
input x_1906;
input x_1907;
input x_1908;
input x_1909;
input x_1910;
input x_1911;
input x_1912;
input x_1913;
input x_1914;
input x_1915;
input x_1916;
input x_1917;
input x_1918;
input x_1919;
input x_1920;
input x_1921;
input x_1922;
input x_1923;
input x_1924;
input x_1925;
input x_1926;
input x_1927;
input x_1928;
input x_1929;
input x_1930;
input x_1931;
input x_1932;
input x_1933;
input x_1934;
input x_1935;
input x_1936;
input x_1937;
input x_1938;
input x_1939;
input x_1940;
input x_1941;
input x_1942;
input x_1943;
input x_1944;
input x_1945;
input x_1946;
input x_1947;
input x_1948;
input x_1949;
input x_1950;
input x_1951;
input x_1952;
input x_1953;
input x_1954;
input x_1955;
input x_1956;
input x_1957;
input x_1958;
input x_1959;
input x_1960;
input x_1961;
input x_1962;
input x_1963;
input x_1964;
input x_1965;
input x_1966;
input x_1967;
input x_1968;
input x_1969;
input x_1970;
input x_1971;
input x_1972;
input x_1973;
input x_1974;
input x_1975;
input x_1976;
input x_1977;
input x_1978;
input x_1979;
input x_1980;
input x_1981;
input x_1982;
input x_1983;
input x_1984;
input x_1985;
input x_1986;
input x_1987;
input x_1988;
input x_1989;
input x_1990;
input x_1991;
input x_1992;
input x_1993;
input x_1994;
input x_1995;
input x_1996;
input x_1997;
input x_1998;
input x_1999;
input x_2000;
input x_2001;
input x_2002;
input x_2003;
input x_2004;
input x_2005;
input x_2006;
input x_2007;
input x_2008;
input x_2009;
input x_2010;
input x_2011;
input x_2012;
input x_2013;
input x_2014;
input x_2015;
input x_2016;
input x_2017;
input x_2018;
input x_2019;
input x_2020;
input x_2021;
input x_2022;
input x_2023;
input x_2024;
input x_2025;
input x_2026;
input x_2027;
input x_2028;
input x_2029;
input x_2030;
input x_2031;
input x_2032;
input x_2033;
input x_2034;
input x_2035;
input x_2036;
input x_2037;
input x_2038;
input x_2039;
input x_2040;
input x_2041;
input x_2042;
input x_2043;
input x_2044;
input x_2045;
input x_2046;
input x_2047;
input x_2048;
input x_2049;
input x_2050;
input x_2051;
input x_2052;
input x_2053;
input x_2054;
input x_2055;
input x_2056;
input x_2057;
input x_2058;
input x_2059;
input x_2060;
input x_2061;
input x_2062;
input x_2063;
input x_2064;
input x_2065;
input x_2066;
input x_2067;
input x_2068;
input x_2069;
input x_2070;
input x_2071;
input x_2072;
input x_2073;
input x_2074;
input x_2075;
input x_2076;
input x_2077;
input x_2078;
input x_2079;
input x_2080;
input x_2081;
input x_2082;
input x_2083;
input x_2084;
input x_2085;
input x_2086;
input x_2087;
input x_2088;
input x_2089;
input x_2090;
input x_2091;
input x_2092;
input x_2093;
input x_2094;
input x_2095;
input x_2096;
input x_2097;
input x_2098;
input x_2099;
input x_2100;
input x_2101;
input x_2102;
input x_2103;
input x_2104;
input x_2105;
input x_2106;
input x_2107;
input x_2108;
input x_2109;
input x_2110;
input x_2111;
input x_2112;
input x_2113;
input x_2114;
input x_2115;
input x_2116;
input x_2117;
input x_2118;
input x_2119;
input x_2120;
input x_2121;
input x_2122;
input x_2123;
input x_2124;
input x_2125;
input x_2126;
input x_2127;
input x_2128;
input x_2129;
input x_2130;
input x_2131;
input x_2132;
input x_2133;
input x_2134;
input x_2135;
input x_2136;
input x_2137;
input x_2138;
input x_2139;
input x_2140;
input x_2141;
input x_2142;
input x_2143;
input x_2144;
input x_2145;
input x_2146;
input x_2147;
input x_2148;
input x_2149;
input x_2150;
input x_2151;
input x_2152;
input x_2153;
input x_2154;
input x_2155;
input x_2156;
input x_2157;
input x_2158;
input x_2159;
input x_2160;
input x_2161;
input x_2162;
input x_2163;
input x_2164;
input x_2165;
input x_2166;
input x_2167;
input x_2168;
input x_2169;
input x_2170;
input x_2171;
input x_2172;
input x_2173;
input x_2174;
input x_2175;
input x_2176;
input x_2177;
input x_2178;
input x_2179;
input x_2180;
input x_2181;
input x_2182;
input x_2183;
input x_2184;
input x_2185;
input x_2186;
input x_2187;
input x_2188;
input x_2189;
input x_2190;
input x_2191;
input x_2192;
input x_2193;
input x_2194;
input x_2195;
input x_2196;
input x_2197;
input x_2198;
input x_2199;
input x_2200;
input x_2201;
input x_2202;
input x_2203;
input x_2204;
input x_2205;
input x_2206;
input x_2207;
input x_2208;
input x_2209;
input x_2210;
input x_2211;
input x_2212;
input x_2213;
input x_2214;
input x_2215;
input x_2216;
input x_2217;
input x_2218;
input x_2219;
input x_2220;
input x_2221;
input x_2222;
input x_2223;
input x_2224;
input x_2225;
input x_2226;
input x_2227;
input x_2228;
input x_2229;
input x_2230;
input x_2231;
input x_2232;
input x_2233;
input x_2234;
input x_2235;
input x_2236;
input x_2237;
input x_2238;
input x_2239;
input x_2240;
input x_2241;
input x_2242;
input x_2243;
input x_2244;
input x_2245;
input x_2246;
input x_2247;
input x_2248;
input x_2249;
input x_2250;
input x_2251;
input x_2252;
input x_2253;
input x_2254;
input x_2255;
input x_2256;
input x_2257;
input x_2258;
input x_2259;
input x_2260;
input x_2261;
input x_2262;
input x_2263;
input x_2264;
input x_2265;
input x_2266;
input x_2267;
input x_2268;
input x_2269;
input x_2270;
input x_2271;
input x_2272;
input x_2273;
input x_2274;
input x_2275;
input x_2276;
input x_2277;
input x_2278;
input x_2279;
input x_2280;
input x_2281;
input x_2282;
input x_2283;
input x_2284;
input x_2285;
input x_2286;
input x_2287;
input x_2288;
input x_2289;
input x_2290;
input x_2291;
input x_2292;
input x_2293;
input x_2294;
input x_2295;
input x_2296;
input x_2297;
input x_2298;
input x_2299;
input x_2300;
input x_2301;
input x_2302;
input x_2303;
input x_2304;
input x_2305;
input x_2306;
input x_2307;
input x_2308;
input x_2309;
input x_2310;
input x_2311;
input x_2312;
input x_2313;
input x_2314;
input x_2315;
input x_2316;
input x_2317;
input x_2318;
input x_2319;
input x_2320;
input x_2321;
input x_2322;
input x_2323;
input x_2324;
input x_2325;
input x_2326;
input x_2327;
input x_2328;
input x_2329;
input x_2330;
input x_2331;
input x_2332;
input x_2333;
input x_2334;
input x_2335;
input x_2336;
input x_2337;
input x_2338;
input x_2339;
input x_2340;
input x_2341;
input x_2342;
input x_2343;
input x_2344;
input x_2345;
input x_2346;
input x_2347;
input x_2348;
input x_2349;
input x_2350;
input x_2351;
input x_2352;
input x_2353;
input x_2354;
input x_2355;
input x_2356;
input x_2357;
input x_2358;
input x_2359;
input x_2360;
input x_2361;
input x_2362;
input x_2363;
input x_2364;
input x_2365;
input x_2366;
input x_2367;
input x_2368;
input x_2369;
input x_2370;
input x_2371;
input x_2372;
input x_2373;
input x_2374;
input x_2375;
input x_2376;
input x_2377;
input x_2378;
input x_2379;
input x_2380;
input x_2381;
input x_2382;
input x_2383;
input x_2384;
input x_2385;
input x_2386;
input x_2387;
input x_2388;
input x_2389;
input x_2390;
input x_2391;
input x_2392;
input x_2393;
input x_2394;
input x_2395;
input x_2396;
input x_2397;
input x_2398;
input x_2399;
input x_2400;
input x_2401;
input x_2402;
input x_2403;
input x_2404;
input x_2405;
input x_2406;
input x_2407;
input x_2408;
input x_2409;
input x_2410;
input x_2411;
input x_2412;
input x_2413;
input x_2414;
input x_2415;
input x_2416;
input x_2417;
input x_2418;
input x_2419;
input x_2420;
input x_2421;
input x_2422;
input x_2423;
input x_2424;
input x_2425;
input x_2426;
input x_2427;
input x_2428;
input x_2429;
input x_2430;
input x_2431;
input x_2432;
input x_2433;
input x_2434;
input x_2435;
input x_2436;
input x_2437;
input x_2438;
input x_2439;
input x_2440;
input x_2441;
input x_2442;
input x_2443;
input x_2444;
input x_2445;
input x_2446;
input x_2447;
input x_2448;
input x_2449;
input x_2450;
input x_2451;
input x_2452;
input x_2453;
input x_2454;
input x_2455;
input x_2456;
input x_2457;
input x_2458;
input x_2459;
input x_2460;
input x_2461;
input x_2462;
input x_2463;
input x_2464;
input x_2465;
input x_2466;
input x_2467;
input x_2468;
input x_2469;
input x_2470;
input x_2471;
input x_2472;
input x_2473;
input x_2474;
input x_2475;
input x_2476;
input x_2477;
input x_2478;
input x_2479;
input x_2480;
input x_2481;
input x_2482;
input x_2483;
input x_2484;
input x_2485;
input x_2486;
input x_2487;
input x_2488;
input x_2489;
input x_2490;
input x_2491;
input x_2492;
input x_2493;
input x_2494;
input x_2495;
input x_2496;
input x_2497;
input x_2498;
input x_2499;
input x_2500;
input x_2501;
input x_2502;
input x_2503;
input x_2504;
input x_2505;
input x_2506;
input x_2507;
input x_2508;
input x_2509;
input x_2510;
input x_2511;
input x_2512;
input x_2513;
input x_2514;
input x_2515;
input x_2516;
input x_2517;
input x_2518;
input x_2519;
input x_2520;
input x_2521;
input x_2522;
input x_2523;
input x_2524;
input x_2525;
input x_2526;
input x_2527;
input x_2528;
input x_2529;
input x_2530;
input x_2531;
input x_2532;
input x_2533;
input x_2534;
input x_2535;
input x_2536;
input x_2537;
input x_2538;
input x_2539;
input x_2540;
input x_2541;
input x_2542;
input x_2543;
input x_2544;
input x_2545;
input x_2546;
input x_2547;
input x_2548;
input x_2549;
input x_2550;
input x_2551;
input x_2552;
input x_2553;
input x_2554;
input x_2555;
input x_2556;
input x_2557;
input x_2558;
input x_2559;
input x_2560;
input x_2561;
input x_2562;
input x_2563;
input x_2564;
input x_2565;
input x_2566;
input x_2567;
input x_2568;
input x_2569;
input x_2570;
input x_2571;
input x_2572;
input x_2573;
input x_2574;
input x_2575;
input x_2576;
input x_2577;
input x_2578;
input x_2579;
input x_2580;
input x_2581;
input x_2582;
input x_2583;
input x_2584;
input x_2585;
input x_2586;
input x_2587;
input x_2588;
input x_2589;
input x_2590;
input x_2591;
input x_2592;
input x_2593;
input x_2594;
input x_2595;
input x_2596;
input x_2597;
input x_2598;
input x_2599;
input x_2600;
input x_2601;
input x_2602;
input x_2603;
input x_2604;
input x_2605;
input x_2606;
input x_2607;
input x_2608;
input x_2609;
input x_2610;
input x_2611;
input x_2612;
input x_2613;
input x_2614;
input x_2615;
input x_2616;
input x_2617;
input x_2618;
input x_2619;
input x_2620;
input x_2621;
input x_2622;
input x_2623;
input x_2624;
input x_2625;
input x_2626;
input x_2627;
input x_2628;
input x_2629;
input x_2630;
input x_2631;
input x_2632;
input x_2633;
input x_2634;
input x_2635;
input x_2636;
input x_2637;
input x_2638;
input x_2639;
input x_2640;
input x_2641;
input x_2642;
input x_2643;
input x_2644;
input x_2645;
input x_2646;
input x_2647;
input x_2648;
input x_2649;
input x_2650;
input x_2651;
input x_2652;
input x_2653;
input x_2654;
input x_2655;
input x_2656;
input x_2657;
input x_2658;
input x_2659;
input x_2660;
input x_2661;
input x_2662;
input x_2663;
input x_2664;
input x_2665;
input x_2666;
input x_2667;
input x_2668;
input x_2669;
input x_2670;
input x_2671;
input x_2672;
input x_2673;
input x_2674;
input x_2675;
input x_2676;
input x_2677;
input x_2678;
input x_2679;
input x_2680;
input x_2681;
input x_2682;
input x_2683;
input x_2684;
input x_2685;
input x_2686;
input x_2687;
input x_2688;
input x_2689;
input x_2690;
input x_2691;
input x_2692;
input x_2693;
input x_2694;
input x_2695;
input x_2696;
input x_2697;
input x_2698;
input x_2699;
input x_2700;
input x_2701;
input x_2702;
input x_2703;
input x_2704;
input x_2705;
input x_2706;
input x_2707;
input x_2708;
input x_2709;
input x_2710;
input x_2711;
input x_2712;
input x_2713;
input x_2714;
input x_2715;
input x_2716;
input x_2717;
input x_2718;
input x_2719;
input x_2720;
input x_2721;
input x_2722;
input x_2723;
input x_2724;
input x_2725;
input x_2726;
input x_2727;
input x_2728;
input x_2729;
input x_2730;
input x_2731;
input x_2732;
input x_2733;
input x_2734;
input x_2735;
input x_2736;
input x_2737;
input x_2738;
input x_2739;
input x_2740;
input x_2741;
input x_2742;
input x_2743;
input x_2744;
input x_2745;
input x_2746;
input x_2747;
input x_2748;
input x_2749;
input x_2750;
input x_2751;
input x_2752;
input x_2753;
input x_2754;
input x_2755;
input x_2756;
input x_2757;
input x_2758;
input x_2759;
input x_2760;
input x_2761;
input x_2762;
input x_2763;
input x_2764;
input x_2765;
input x_2766;
input x_2767;
input x_2768;
input x_2769;
input x_2770;
input x_2771;
input x_2772;
input x_2773;
input x_2774;
input x_2775;
input x_2776;
input x_2777;
input x_2778;
input x_2779;
input x_2780;
input x_2781;
input x_2782;
input x_2783;
input x_2784;
input x_2785;
input x_2786;
input x_2787;
input x_2788;
input x_2789;
input x_2790;
input x_2791;
input x_2792;
input x_2793;
input x_2794;
input x_2795;
input x_2796;
input x_2797;
input x_2798;
input x_2799;
input x_2800;
input x_2801;
input x_2802;
input x_2803;
input x_2804;
input x_2805;
input x_2806;
input x_2807;
input x_2808;
input x_2809;
input x_2810;
input x_2811;
input x_2812;
input x_2813;
input x_2814;
input x_2815;
input x_2816;
input x_2817;
input x_2818;
input x_2819;
input x_2820;
input x_2821;
input x_2822;
input x_2823;
input x_2824;
input x_2825;
input x_2826;
input x_2827;
input x_2828;
input x_2829;
input x_2830;
input x_2831;
input x_2832;
input x_2833;
input x_2834;
input x_2835;
input x_2836;
input x_2837;
input x_2838;
input x_2839;
input x_2840;
input x_2841;
input x_2842;
input x_2843;
input x_2844;
input x_2845;
input x_2846;
input x_2847;
input x_2848;
input x_2849;
input x_2850;
input x_2851;
input x_2852;
input x_2853;
input x_2854;
input x_2855;
input x_2856;
input x_2857;
input x_2858;
input x_2859;
input x_2860;
input x_2861;
input x_2862;
input x_2863;
input x_2864;
input x_2865;
input x_2866;
input x_2867;
input x_2868;
input x_2869;
input x_2870;
input x_2871;
input x_2872;
input x_2873;
input x_2874;
input x_2875;
input x_2876;
input x_2877;
input x_2878;
input x_2879;
input x_2880;
input x_2881;
input x_2882;
input x_2883;
input x_2884;
input x_2885;
input x_2886;
input x_2887;
input x_2888;
input x_2889;
input x_2890;
input x_2891;
input x_2892;
input x_2893;
input x_2894;
input x_2895;
input x_2896;
input x_2897;
input x_2898;
input x_2899;
input x_2900;
input x_2901;
input x_2902;
input x_2903;
input x_2904;
input x_2905;
input x_2906;
input x_2907;
input x_2908;
input x_2909;
input x_2910;
input x_2911;
input x_2912;
input x_2913;
input x_2914;
input x_2915;
input x_2916;
input x_2917;
input x_2918;
input x_2919;
input x_2920;
input x_2921;
input x_2922;
input x_2923;
input x_2924;
input x_2925;
input x_2926;
input x_2927;
input x_2928;
input x_2929;
input x_2930;
input x_2931;
input x_2932;
input x_2933;
input x_2934;
input x_2935;
input x_2936;
input x_2937;
input x_2938;
input x_2939;
input x_2940;
input x_2941;
input x_2942;
input x_2943;
input x_2944;
input x_2945;
input x_2946;
input x_2947;
input x_2948;
input x_2949;
input x_2950;
input x_2951;
input x_2952;
input x_2953;
input x_2954;
input x_2955;
input x_2956;
input x_2957;
input x_2958;
input x_2959;
input x_2960;
input x_2961;
input x_2962;
input x_2963;
input x_2964;
input x_2965;
input x_2966;
input x_2967;
input x_2968;
input x_2969;
input x_2970;
input x_2971;
input x_2972;
input x_2973;
input x_2974;
input x_2975;
input x_2976;
input x_2977;
input x_2978;
input x_2979;
input x_2980;
input x_2981;
input x_2982;
input x_2983;
input x_2984;
input x_2985;
input x_2986;
input x_2987;
input x_2988;
input x_2989;
input x_2990;
input x_2991;
input x_2992;
input x_2993;
input x_2994;
input x_2995;
input x_2996;
input x_2997;
input x_2998;
input x_2999;
input x_3000;
input x_3001;
input x_3002;
input x_3003;
input x_3004;
input x_3005;
input x_3006;
input x_3007;
input x_3008;
input x_3009;
input x_3010;
input x_3011;
input x_3012;
input x_3013;
input x_3014;
input x_3015;
input x_3016;
input x_3017;
input x_3018;
input x_3019;
input x_3020;
input x_3021;
input x_3022;
input x_3023;
input x_3024;
input x_3025;
input x_3026;
input x_3027;
input x_3028;
input x_3029;
input x_3030;
input x_3031;
input x_3032;
input x_3033;
input x_3034;
input x_3035;
input x_3036;
input x_3037;
input x_3038;
input x_3039;
input x_3040;
input x_3041;
input x_3042;
input x_3043;
input x_3044;
input x_3045;
input x_3046;
input x_3047;
input x_3048;
input x_3049;
input x_3050;
input x_3051;
input x_3052;
input x_3053;
input x_3054;
input x_3055;
input x_3056;
input x_3057;
input x_3058;
input x_3059;
input x_3060;
input x_3061;
input x_3062;
input x_3063;
input x_3064;
input x_3065;
input x_3066;
input x_3067;
input x_3068;
input x_3069;
input x_3070;
input x_3071;
input x_3072;
input x_3073;
input x_3074;
input x_3075;
input x_3076;
input x_3077;
input x_3078;
input x_3079;
input x_3080;
input x_3081;
input x_3082;
input x_3083;
input x_3084;
input x_3085;
input x_3086;
input x_3087;
input x_3088;
input x_3089;
input x_3090;
input x_3091;
input x_3092;
input x_3093;
input x_3094;
input x_3095;
input x_3096;
input x_3097;
input x_3098;
input x_3099;
input x_3100;
input x_3101;
input x_3102;
input x_3103;
input x_3104;
input x_3105;
input x_3106;
input x_3107;
input x_3108;
input x_3109;
input x_3110;
input x_3111;
input x_3112;
input x_3113;
input x_3114;
input x_3115;
input x_3116;
input x_3117;
input x_3118;
input x_3119;
input x_3120;
input x_3121;
input x_3122;
input x_3123;
input x_3124;
input x_3125;
input x_3126;
input x_3127;
input x_3128;
input x_3129;
input x_3130;
input x_3131;
input x_3132;
input x_3133;
input x_3134;
input x_3135;
input x_3136;
input x_3137;
input x_3138;
input x_3139;
input x_3140;
input x_3141;
input x_3142;
input x_3143;
input x_3144;
input x_3145;
input x_3146;
input x_3147;
input x_3148;
input x_3149;
input x_3150;
input x_3151;
input x_3152;
input x_3153;
input x_3154;
input x_3155;
input x_3156;
input x_3157;
input x_3158;
input x_3159;
input x_3160;
input x_3161;
input x_3162;
input x_3163;
input x_3164;
input x_3165;
input x_3166;
input x_3167;
input x_3168;
input x_3169;
input x_3170;
input x_3171;
input x_3172;
input x_3173;
input x_3174;
input x_3175;
input x_3176;
input x_3177;
input x_3178;
input x_3179;
input x_3180;
input x_3181;
input x_3182;
input x_3183;
input x_3184;
input x_3185;
input x_3186;
input x_3187;
input x_3188;
input x_3189;
input x_3190;
input x_3191;
input x_3192;
input x_3193;
input x_3194;
input x_3195;
input x_3196;
input x_3197;
input x_3198;
input x_3199;
input x_3200;
input x_3201;
input x_3202;
input x_3203;
input x_3204;
input x_3205;
input x_3206;
input x_3207;
input x_3208;
input x_3209;
input x_3210;
input x_3211;
input x_3212;
input x_3213;
input x_3214;
input x_3215;
input x_3216;
input x_3217;
input x_3218;
input x_3219;
input x_3220;
input x_3221;
input x_3222;
input x_3223;
input x_3224;
input x_3225;
input x_3226;
input x_3227;
input x_3228;
input x_3229;
input x_3230;
input x_3231;
input x_3232;
input x_3233;
input x_3234;
input x_3235;
input x_3236;
input x_3237;
input x_3238;
input x_3239;
input x_3240;
input x_3241;
input x_3242;
input x_3243;
input x_3244;
input x_3245;
input x_3246;
input x_3247;
input x_3248;
input x_3249;
input x_3250;
input x_3251;
input x_3252;
input x_3253;
input x_3254;
input x_3255;
input x_3256;
input x_3257;
input x_3258;
input x_3259;
input x_3260;
input x_3261;
input x_3262;
input x_3263;
input x_3264;
input x_3265;
input x_3266;
input x_3267;
input x_3268;
input x_3269;
input x_3270;
input x_3271;
input x_3272;
input x_3273;
input x_3274;
input x_3275;
input x_3276;
input x_3277;
input x_3278;
input x_3279;
input x_3280;
input x_3281;
input x_3282;
input x_3283;
input x_3284;
input x_3285;
input x_3286;
input x_3287;
input x_3288;
input x_3289;
input x_3290;
input x_3291;
input x_3292;
input x_3293;
input x_3294;
input x_3295;
input x_3296;
input x_3297;
input x_3298;
input x_3299;
input x_3300;
input x_3301;
input x_3302;
input x_3303;
input x_3304;
input x_3305;
input x_3306;
input x_3307;
input x_3308;
input x_3309;
input x_3310;
input x_3311;
input x_3312;
input x_3313;
input x_3314;
input x_3315;
input x_3316;
input x_3317;
input x_3318;
input x_3319;
input x_3320;
input x_3321;
input x_3322;
input x_3323;
input x_3324;
input x_3325;
input x_3326;
input x_3327;
input x_3328;
input x_3329;
input x_3330;
input x_3331;
input x_3332;
input x_3333;
input x_3334;
input x_3335;
input x_3336;
input x_3337;
input x_3338;
input x_3339;
input x_3340;
input x_3341;
input x_3342;
input x_3343;
input x_3344;
input x_3345;
input x_3346;
input x_3347;
input x_3348;
input x_3349;
input x_3350;
input x_3351;
input x_3352;
input x_3353;
input x_3354;
input x_3355;
input x_3356;
input x_3357;
input x_3358;
input x_3359;
input x_3360;
input x_3361;
input x_3362;
input x_3363;
input x_3364;
input x_3365;
input x_3366;
input x_3367;
input x_3368;
input x_3369;
input x_3370;
input x_3371;
input x_3372;
input x_3373;
input x_3374;
input x_3375;
input x_3376;
input x_3377;
input x_3378;
input x_3379;
input x_3380;
input x_3381;
input x_3382;
input x_3383;
input x_3384;
input x_3385;
input x_3386;
input x_3387;
input x_3388;
input x_3389;
input x_3390;
input x_3391;
input x_3392;
input x_3393;
input x_3394;
input x_3395;
input x_3396;
input x_3397;
input x_3398;
input x_3399;
input x_3400;
input x_3401;
input x_3402;
input x_3403;
input x_3404;
input x_3405;
input x_3406;
input x_3407;
input x_3408;
input x_3409;
input x_3410;
input x_3411;
input x_3412;
input x_3413;
input x_3414;
input x_3415;
input x_3416;
input x_3417;
input x_3418;
input x_3419;
input x_3420;
input x_3421;
input x_3422;
input x_3423;
input x_3424;
input x_3425;
input x_3426;
input x_3427;
input x_3428;
input x_3429;
input x_3430;
input x_3431;
input x_3432;
input x_3433;
input x_3434;
input x_3435;
input x_3436;
input x_3437;
input x_3438;
input x_3439;
input x_3440;
input x_3441;
input x_3442;
input x_3443;
input x_3444;
input x_3445;
input x_3446;
input x_3447;
input x_3448;
input x_3449;
input x_3450;
input x_3451;
input x_3452;
input x_3453;
input x_3454;
input x_3455;
input x_3456;
input x_3457;
input x_3458;
input x_3459;
input x_3460;
input x_3461;
input x_3462;
input x_3463;
input x_3464;
input x_3465;
input x_3466;
input x_3467;
input x_3468;
input x_3469;
input x_3470;
input x_3471;
input x_3472;
input x_3473;
input x_3474;
input x_3475;
input x_3476;
input x_3477;
input x_3478;
input x_3479;
input x_3480;
input x_3481;
input x_3482;
input x_3483;
input x_3484;
input x_3485;
input x_3486;
input x_3487;
input x_3488;
input x_3489;
input x_3490;
input x_3491;
input x_3492;
input x_3493;
input x_3494;
input x_3495;
input x_3496;
input x_3497;
input x_3498;
input x_3499;
input x_3500;
input x_3501;
input x_3502;
input x_3503;
input x_3504;
input x_3505;
input x_3506;
input x_3507;
input x_3508;
input x_3509;
input x_3510;
input x_3511;
input x_3512;
input x_3513;
input x_3514;
input x_3515;
input x_3516;
input x_3517;
input x_3518;
input x_3519;
input x_3520;
input x_3521;
input x_3522;
input x_3523;
input x_3524;
input x_3525;
input x_3526;
input x_3527;
input x_3528;
input x_3529;
input x_3530;
input x_3531;
input x_3532;
input x_3533;
input x_3534;
input x_3535;
input x_3536;
input x_3537;
input x_3538;
input x_3539;
input x_3540;
input x_3541;
input x_3542;
input x_3543;
input x_3544;
input x_3545;
input x_3546;
input x_3547;
input x_3548;
input x_3549;
input x_3550;
input x_3551;
input x_3552;
input x_3553;
input x_3554;
input x_3555;
input x_3556;
input x_3557;
input x_3558;
input x_3559;
input x_3560;
input x_3561;
input x_3562;
input x_3563;
input x_3564;
input x_3565;
input x_3566;
input x_3567;
input x_3568;
input x_3569;
input x_3570;
input x_3571;
input x_3572;
input x_3573;
input x_3574;
input x_3575;
input x_3576;
input x_3577;
input x_3578;
input x_3579;
input x_3580;
input x_3581;
input x_3582;
input x_3583;
input x_3584;
input x_3585;
input x_3586;
input x_3587;
input x_3588;
input x_3589;
input x_3590;
input x_3591;
input x_3592;
input x_3593;
input x_3594;
input x_3595;
input x_3596;
input x_3597;
input x_3598;
input x_3599;
input x_3600;
input x_3601;
input x_3602;
input x_3603;
input x_3604;
input x_3605;
input x_3606;
input x_3607;
input x_3608;
input x_3609;
input x_3610;
input x_3611;
input x_3612;
input x_3613;
input x_3614;
input x_3615;
input x_3616;
input x_3617;
input x_3618;
input x_3619;
input x_3620;
input x_3621;
input x_3622;
input x_3623;
input x_3624;
input x_3625;
input x_3626;
input x_3627;
input x_3628;
input x_3629;
input x_3630;
input x_3631;
input x_3632;
input x_3633;
input x_3634;
input x_3635;
input x_3636;
input x_3637;
input x_3638;
input x_3639;
input x_3640;
input x_3641;
input x_3642;
input x_3643;
input x_3644;
input x_3645;
input x_3646;
input x_3647;
input x_3648;
input x_3649;
input x_3650;
input x_3651;
input x_3652;
input x_3653;
input x_3654;
input x_3655;
input x_3656;
input x_3657;
input x_3658;
input x_3659;
input x_3660;
input x_3661;
input x_3662;
input x_3663;
input x_3664;
input x_3665;
input x_3666;
input x_3667;
input x_3668;
input x_3669;
input x_3670;
input x_3671;
input x_3672;
input x_3673;
input x_3674;
input x_3675;
input x_3676;
input x_3677;
input x_3678;
input x_3679;
input x_3680;
input x_3681;
input x_3682;
input x_3683;
input x_3684;
input x_3685;
input x_3686;
input x_3687;
input x_3688;
input x_3689;
input x_3690;
input x_3691;
input x_3692;
input x_3693;
input x_3694;
input x_3695;
input x_3696;
input x_3697;
input x_3698;
input x_3699;
input x_3700;
input x_3701;
input x_3702;
input x_3703;
input x_3704;
input x_3705;
input x_3706;
input x_3707;
input x_3708;
input x_3709;
input x_3710;
input x_3711;
input x_3712;
input x_3713;
input x_3714;
input x_3715;
input x_3716;
input x_3717;
input x_3718;
input x_3719;
input x_3720;
input x_3721;
input x_3722;
input x_3723;
input x_3724;
input x_3725;
input x_3726;
input x_3727;
input x_3728;
input x_3729;
input x_3730;
input x_3731;
input x_3732;
input x_3733;
input x_3734;
input x_3735;
input x_3736;
input x_3737;
input x_3738;
input x_3739;
input x_3740;
input x_3741;
input x_3742;
input x_3743;
input x_3744;
input x_3745;
input x_3746;
input x_3747;
input x_3748;
input x_3749;
input x_3750;
input x_3751;
input x_3752;
input x_3753;
input x_3754;
input x_3755;
input x_3756;
input x_3757;
input x_3758;
input x_3759;
input x_3760;
input x_3761;
input x_3762;
input x_3763;
input x_3764;
input x_3765;
input x_3766;
input x_3767;
input x_3768;
input x_3769;
input x_3770;
input x_3771;
input x_3772;
input x_3773;
input x_3774;
input x_3775;
input x_3776;
input x_3777;
input x_3778;
input x_3779;
input x_3780;
input x_3781;
input x_3782;
input x_3783;
input x_3784;
input x_3785;
input x_3786;
input x_3787;
input x_3788;
input x_3789;
input x_3790;
input x_3791;
input x_3792;
input x_3793;
input x_3794;
input x_3795;
input x_3796;
input x_3797;
input x_3798;
input x_3799;
input x_3800;
input x_3801;
input x_3802;
input x_3803;
input x_3804;
input x_3805;
input x_3806;
input x_3807;
input x_3808;
input x_3809;
input x_3810;
input x_3811;
input x_3812;
input x_3813;
input x_3814;
input x_3815;
input x_3816;
input x_3817;
input x_3818;
input x_3819;
input x_3820;
input x_3821;
input x_3822;
input x_3823;
input x_3824;
input x_3825;
input x_3826;
input x_3827;
input x_3828;
input x_3829;
input x_3830;
input x_3831;
input x_3832;
input x_3833;
input x_3834;
input x_3835;
input x_3836;
input x_3837;
input x_3838;
input x_3839;
input x_3840;
input x_3841;
input x_3842;
input x_3843;
input x_3844;
input x_3845;
input x_3846;
input x_3847;
input x_3848;
input x_3849;
input x_3850;
input x_3851;
input x_3852;
input x_3853;
input x_3854;
input x_3855;
input x_3856;
input x_3857;
input x_3858;
input x_3859;
input x_3860;
input x_3861;
input x_3862;
input x_3863;
input x_3864;
input x_3865;
input x_3866;
input x_3867;
input x_3868;
input x_3869;
input x_3870;
input x_3871;
input x_3872;
input x_3873;
input x_3874;
input x_3875;
input x_3876;
input x_3877;
input x_3878;
input x_3879;
input x_3880;
input x_3881;
input x_3882;
input x_3883;
input x_3884;
input x_3885;
input x_3886;
input x_3887;
input x_3888;
input x_3889;
input x_3890;
input x_3891;
input x_3892;
input x_3893;
input x_3894;
input x_3895;
input x_3896;
input x_3897;
input x_3898;
input x_3899;
input x_3900;
input x_3901;
input x_3902;
input x_3903;
input x_3904;
input x_3905;
input x_3906;
input x_3907;
input x_3908;
input x_3909;
input x_3910;
input x_3911;
input x_3912;
input x_3913;
input x_3914;
input x_3915;
input x_3916;
input x_3917;
input x_3918;
input x_3919;
input x_3920;
input x_3921;
input x_3922;
input x_3923;
input x_3924;
input x_3925;
input x_3926;
input x_3927;
input x_3928;
input x_3929;
input x_3930;
input x_3931;
input x_3932;
input x_3933;
input x_3934;
input x_3935;
input x_3936;
input x_3937;
input x_3938;
input x_3939;
input x_3940;
input x_3941;
input x_3942;
input x_3943;
input x_3944;
input x_3945;
input x_3946;
input x_3947;
input x_3948;
input x_3949;
input x_3950;
input x_3951;
input x_3952;
input x_3953;
input x_3954;
input x_3955;
input x_3956;
input x_3957;
input x_3958;
input x_3959;
input x_3960;
input x_3961;
input x_3962;
input x_3963;
input x_3964;
input x_3965;
input x_3966;
input x_3967;
input x_3968;
input x_3969;
input x_3970;
input x_3971;
input x_3972;
input x_3973;
input x_3974;
input x_3975;
input x_3976;
input x_3977;
input x_3978;
input x_3979;
input x_3980;
input x_3981;
input x_3982;
input x_3983;
input x_3984;
input x_3985;
input x_3986;
input x_3987;
input x_3988;
input x_3989;
input x_3990;
input x_3991;
input x_3992;
input x_3993;
input x_3994;
input x_3995;
input x_3996;
input x_3997;
input x_3998;
input x_3999;
input x_4000;
input x_4001;
input x_4002;
input x_4003;
input x_4004;
input x_4005;
input x_4006;
input x_4007;
input x_4008;
input x_4009;
input x_4010;
input x_4011;
input x_4012;
input x_4013;
input x_4014;
input x_4015;
input x_4016;
input x_4017;
input x_4018;
input x_4019;
input x_4020;
input x_4021;
input x_4022;
input x_4023;
input x_4024;
input x_4025;
input x_4026;
input x_4027;
input x_4028;
input x_4029;
input x_4030;
input x_4031;
input x_4032;
input x_4033;
input x_4034;
input x_4035;
input x_4036;
input x_4037;
input x_4038;
input x_4039;
input x_4040;
input x_4041;
input x_4042;
input x_4043;
input x_4044;
input x_4045;
input x_4046;
input x_4047;
input x_4048;
input x_4049;
input x_4050;
input x_4051;
input x_4052;
input x_4053;
input x_4054;
input x_4055;
input x_4056;
input x_4057;
input x_4058;
input x_4059;
input x_4060;
input x_4061;
input x_4062;
input x_4063;
input x_4064;
input x_4065;
input x_4066;
input x_4067;
input x_4068;
input x_4069;
input x_4070;
input x_4071;
input x_4072;
input x_4073;
input x_4074;
input x_4075;
input x_4076;
input x_4077;
input x_4078;
input x_4079;
input x_4080;
input x_4081;
input x_4082;
input x_4083;
input x_4084;
input x_4085;
input x_4086;
input x_4087;
input x_4088;
input x_4089;
input x_4090;
input x_4091;
input x_4092;
input x_4093;
input x_4094;
input x_4095;
input x_4096;
input x_4097;
input x_4098;
input x_4099;
input x_4100;
input x_4101;
input x_4102;
input x_4103;
input x_4104;
input x_4105;
input x_4106;
input x_4107;
input x_4108;
input x_4109;
input x_4110;
input x_4111;
input x_4112;
input x_4113;
input x_4114;
input x_4115;
input x_4116;
input x_4117;
input x_4118;
input x_4119;
input x_4120;
input x_4121;
input x_4122;
input x_4123;
input x_4124;
input x_4125;
input x_4126;
input x_4127;
input x_4128;
input x_4129;
input x_4130;
input x_4131;
input x_4132;
input x_4133;
input x_4134;
input x_4135;
input x_4136;
input x_4137;
input x_4138;
input x_4139;
input x_4140;
input x_4141;
input x_4142;
input x_4143;
input x_4144;
input x_4145;
input x_4146;
input x_4147;
input x_4148;
input x_4149;
input x_4150;
input x_4151;
input x_4152;
input x_4153;
input x_4154;
input x_4155;
input x_4156;
input x_4157;
input x_4158;
input x_4159;
input x_4160;
input x_4161;
input x_4162;
input x_4163;
input x_4164;
input x_4165;
input x_4166;
input x_4167;
input x_4168;
input x_4169;
input x_4170;
input x_4171;
input x_4172;
input x_4173;
input x_4174;
input x_4175;
input x_4176;
input x_4177;
input x_4178;
input x_4179;
input x_4180;
input x_4181;
input x_4182;
input x_4183;
input x_4184;
input x_4185;
input x_4186;
input x_4187;
input x_4188;
input x_4189;
input x_4190;
input x_4191;
input x_4192;
input x_4193;
input x_4194;
input x_4195;
input x_4196;
input x_4197;
input x_4198;
input x_4199;
input x_4200;
input x_4201;
input x_4202;
input x_4203;
input x_4204;
input x_4205;
input x_4206;
input x_4207;
input x_4208;
input x_4209;
input x_4210;
input x_4211;
input x_4212;
input x_4213;
input x_4214;
input x_4215;
input x_4216;
input x_4217;
input x_4218;
input x_4219;
input x_4220;
input x_4221;
input x_4222;
input x_4223;
input x_4224;
input x_4225;
input x_4226;
input x_4227;
input x_4228;
input x_4229;
input x_4230;
input x_4231;
input x_4232;
input x_4233;
input x_4234;
input x_4235;
input x_4236;
input x_4237;
input x_4238;
input x_4239;
input x_4240;
input x_4241;
input x_4242;
input x_4243;
input x_4244;
input x_4245;
input x_4246;
input x_4247;
input x_4248;
input x_4249;
input x_4250;
input x_4251;
input x_4252;
input x_4253;
input x_4254;
input x_4255;
input x_4256;
input x_4257;
input x_4258;
input x_4259;
input x_4260;
input x_4261;
input x_4262;
input x_4263;
input x_4264;
input x_4265;
input x_4266;
input x_4267;
input x_4268;
input x_4269;
input x_4270;
input x_4271;
input x_4272;
input x_4273;
input x_4274;
input x_4275;
input x_4276;
input x_4277;
input x_4278;
input x_4279;
input x_4280;
input x_4281;
input x_4282;
input x_4283;
input x_4284;
input x_4285;
input x_4286;
input x_4287;
input x_4288;
input x_4289;
input x_4290;
input x_4291;
input x_4292;
input x_4293;
input x_4294;
input x_4295;
input x_4296;
input x_4297;
input x_4298;
input x_4299;
input x_4300;
input x_4301;
input x_4302;
input x_4303;
input x_4304;
input x_4305;
input x_4306;
input x_4307;
input x_4308;
input x_4309;
input x_4310;
input x_4311;
input x_4312;
input x_4313;
input x_4314;
input x_4315;
input x_4316;
input x_4317;
input x_4318;
input x_4319;
input x_4320;
input x_4321;
input x_4322;
input x_4323;
input x_4324;
input x_4325;
input x_4326;
input x_4327;
input x_4328;
input x_4329;
input x_4330;
input x_4331;
input x_4332;
input x_4333;
input x_4334;
input x_4335;
input x_4336;
input x_4337;
input x_4338;
input x_4339;
input x_4340;
input x_4341;
input x_4342;
input x_4343;
input x_4344;
input x_4345;
input x_4346;
input x_4347;
input x_4348;
input x_4349;
input x_4350;
input x_4351;
input x_4352;
input x_4353;
input x_4354;
input x_4355;
input x_4356;
input x_4357;
input x_4358;
input x_4359;
input x_4360;
input x_4361;
input x_4362;
input x_4363;
input x_4364;
input x_4365;
input x_4366;
input x_4367;
input x_4368;
input x_4369;
input x_4370;
input x_4371;
input x_4372;
input x_4373;
input x_4374;
input x_4375;
input x_4376;
input x_4377;
input x_4378;
input x_4379;
input x_4380;
input x_4381;
input x_4382;
input x_4383;
input x_4384;
input x_4385;
input x_4386;
input x_4387;
input x_4388;
input x_4389;
input x_4390;
input x_4391;
input x_4392;
input x_4393;
input x_4394;
input x_4395;
input x_4396;
input x_4397;
input x_4398;
input x_4399;
input x_4400;
input x_4401;
input x_4402;
input x_4403;
input x_4404;
input x_4405;
input x_4406;
input x_4407;
input x_4408;
input x_4409;
input x_4410;
input x_4411;
input x_4412;
input x_4413;
input x_4414;
input x_4415;
input x_4416;
input x_4417;
input x_4418;
input x_4419;
input x_4420;
input x_4421;
input x_4422;
input x_4423;
input x_4424;
input x_4425;
input x_4426;
input x_4427;
input x_4428;
input x_4429;
input x_4430;
input x_4431;
input x_4432;
input x_4433;
input x_4434;
input x_4435;
input x_4436;
input x_4437;
input x_4438;
input x_4439;
input x_4440;
input x_4441;
input x_4442;
input x_4443;
input x_4444;
input x_4445;
input x_4446;
input x_4447;
input x_4448;
input x_4449;
input x_4450;
input x_4451;
input x_4452;
input x_4453;
input x_4454;
input x_4455;
input x_4456;
input x_4457;
input x_4458;
input x_4459;
input x_4460;
input x_4461;
input x_4462;
input x_4463;
input x_4464;
input x_4465;
input x_4466;
input x_4467;
input x_4468;
input x_4469;
input x_4470;
input x_4471;
input x_4472;
input x_4473;
input x_4474;
input x_4475;
input x_4476;
input x_4477;
input x_4478;
input x_4479;
input x_4480;
input x_4481;
input x_4482;
input x_4483;
input x_4484;
input x_4485;
input x_4486;
input x_4487;
input x_4488;
input x_4489;
input x_4490;
input x_4491;
input x_4492;
input x_4493;
input x_4494;
input x_4495;
input x_4496;
input x_4497;
input x_4498;
input x_4499;
input x_4500;
input x_4501;
input x_4502;
input x_4503;
input x_4504;
input x_4505;
input x_4506;
input x_4507;
input x_4508;
input x_4509;
input x_4510;
input x_4511;
input x_4512;
input x_4513;
input x_4514;
input x_4515;
input x_4516;
input x_4517;
input x_4518;
input x_4519;
input x_4520;
input x_4521;
input x_4522;
input x_4523;
input x_4524;
input x_4525;
input x_4526;
input x_4527;
input x_4528;
input x_4529;
input x_4530;
input x_4531;
input x_4532;
input x_4533;
input x_4534;
input x_4535;
input x_4536;
input x_4537;
input x_4538;
input x_4539;
input x_4540;
input x_4541;
input x_4542;
input x_4543;
input x_4544;
input x_4545;
input x_4546;
input x_4547;
input x_4548;
input x_4549;
input x_4550;
input x_4551;
input x_4552;
input x_4553;
input x_4554;
input x_4555;
input x_4556;
input x_4557;
input x_4558;
input x_4559;
input x_4560;
input x_4561;
input x_4562;
input x_4563;
input x_4564;
input x_4565;
input x_4566;
input x_4567;
input x_4568;
input x_4569;
input x_4570;
input x_4571;
input x_4572;
input x_4573;
input x_4574;
input x_4575;
input x_4576;
input x_4577;
input x_4578;
input x_4579;
input x_4580;
input x_4581;
input x_4582;
input x_4583;
input x_4584;
input x_4585;
input x_4586;
input x_4587;
input x_4588;
input x_4589;
input x_4590;
input x_4591;
input x_4592;
input x_4593;
input x_4594;
input x_4595;
input x_4596;
input x_4597;
input x_4598;
input x_4599;
input x_4600;
input x_4601;
input x_4602;
input x_4603;
input x_4604;
input x_4605;
input x_4606;
input x_4607;
input x_4608;
input x_4609;
input x_4610;
input x_4611;
input x_4612;
input x_4613;
input x_4614;
input x_4615;
input x_4616;
input x_4617;
input x_4618;
input x_4619;
input x_4620;
input x_4621;
input x_4622;
input x_4623;
input x_4624;
input x_4625;
input x_4626;
input x_4627;
input x_4628;
input x_4629;
input x_4630;
input x_4631;
input x_4632;
input x_4633;
input x_4634;
input x_4635;
input x_4636;
input x_4637;
input x_4638;
input x_4639;
input x_4640;
input x_4641;
input x_4642;
input x_4643;
input x_4644;
input x_4645;
input x_4646;
input x_4647;
input x_4648;
input x_4649;
input x_4650;
input x_4651;
input x_4652;
input x_4653;
input x_4654;
input x_4655;
input x_4656;
input x_4657;
input x_4658;
input x_4659;
input x_4660;
input x_4661;
input x_4662;
input x_4663;
input x_4664;
input x_4665;
input x_4666;
input x_4667;
input x_4668;
input x_4669;
input x_4670;
input x_4671;
input x_4672;
input x_4673;
input x_4674;
input x_4675;
input x_4676;
input x_4677;
input x_4678;
input x_4679;
input x_4680;
input x_4681;
input x_4682;
input x_4683;
input x_4684;
input x_4685;
input x_4686;
input x_4687;
input x_4688;
input x_4689;
input x_4690;
input x_4691;
input x_4692;
input x_4693;
input x_4694;
input x_4695;
input x_4696;
input x_4697;
input x_4698;
input x_4699;
input x_4700;
input x_4701;
input x_4702;
input x_4703;
input x_4704;
input x_4705;
input x_4706;
input x_4707;
input x_4708;
input x_4709;
input x_4710;
input x_4711;
input x_4712;
input x_4713;
input x_4714;
input x_4715;
input x_4716;
input x_4717;
input x_4718;
input x_4719;
input x_4720;
input x_4721;
input x_4722;
input x_4723;
input x_4724;
input x_4725;
input x_4726;
input x_4727;
input x_4728;
input x_4729;
input x_4730;
input x_4731;
input x_4732;
input x_4733;
input x_4734;
input x_4735;
input x_4736;
input x_4737;
input x_4738;
input x_4739;
input x_4740;
input x_4741;
input x_4742;
input x_4743;
input x_4744;
input x_4745;
input x_4746;
input x_4747;
input x_4748;
input x_4749;
input x_4750;
input x_4751;
input x_4752;
input x_4753;
input x_4754;
input x_4755;
input x_4756;
input x_4757;
input x_4758;
input x_4759;
input x_4760;
input x_4761;
input x_4762;
input x_4763;
input x_4764;
input x_4765;
input x_4766;
input x_4767;
input x_4768;
input x_4769;
input x_4770;
input x_4771;
input x_4772;
input x_4773;
input x_4774;
input x_4775;
input x_4776;
input x_4777;
input x_4778;
input x_4779;
input x_4780;
input x_4781;
input x_4782;
input x_4783;
input x_4784;
input x_4785;
input x_4786;
input x_4787;
input x_4788;
input x_4789;
input x_4790;
input x_4791;
input x_4792;
input x_4793;
input x_4794;
input x_4795;
input x_4796;
input x_4797;
input x_4798;
input x_4799;
input x_4800;
input x_4801;
input x_4802;
input x_4803;
input x_4804;
input x_4805;
input x_4806;
input x_4807;
input x_4808;
input x_4809;
input x_4810;
input x_4811;
input x_4812;
input x_4813;
input x_4814;
input x_4815;
input x_4816;
input x_4817;
input x_4818;
input x_4819;
input x_4820;
input x_4821;
input x_4822;
input x_4823;
input x_4824;
input x_4825;
input x_4826;
input x_4827;
input x_4828;
input x_4829;
input x_4830;
input x_4831;
input x_4832;
input x_4833;
input x_4834;
input x_4835;
input x_4836;
input x_4837;
input x_4838;
input x_4839;
input x_4840;
input x_4841;
input x_4842;
input x_4843;
input x_4844;
input x_4845;
input x_4846;
input x_4847;
input x_4848;
input x_4849;
input x_4850;
input x_4851;
input x_4852;
input x_4853;
input x_4854;
input x_4855;
input x_4856;
input x_4857;
input x_4858;
input x_4859;
input x_4860;
input x_4861;
input x_4862;
input x_4863;
input x_4864;
input x_4865;
input x_4866;
input x_4867;
input x_4868;
input x_4869;
input x_4870;
input x_4871;
input x_4872;
input x_4873;
input x_4874;
input x_4875;
input x_4876;
input x_4877;
input x_4878;
input x_4879;
input x_4880;
input x_4881;
input x_4882;
input x_4883;
input x_4884;
input x_4885;
input x_4886;
input x_4887;
input x_4888;
input x_4889;
input x_4890;
input x_4891;
input x_4892;
input x_4893;
input x_4894;
input x_4895;
input x_4896;
input x_4897;
input x_4898;
input x_4899;
input x_4900;
input x_4901;
input x_4902;
input x_4903;
input x_4904;
input x_4905;
input x_4906;
input x_4907;
input x_4908;
input x_4909;
input x_4910;
input x_4911;
input x_4912;
input x_4913;
input x_4914;
input x_4915;
input x_4916;
input x_4917;
input x_4918;
input x_4919;
input x_4920;
input x_4921;
input x_4922;
input x_4923;
input x_4924;
input x_4925;
input x_4926;
input x_4927;
input x_4928;
input x_4929;
input x_4930;
input x_4931;
input x_4932;
input x_4933;
input x_4934;
input x_4935;
input x_4936;
input x_4937;
input x_4938;
input x_4939;
input x_4940;
input x_4941;
input x_4942;
input x_4943;
input x_4944;
input x_4945;
input x_4946;
input x_4947;
input x_4948;
input x_4949;
input x_4950;
input x_4951;
input x_4952;
input x_4953;
input x_4954;
input x_4955;
input x_4956;
input x_4957;
input x_4958;
input x_4959;
input x_4960;
input x_4961;
input x_4962;
input x_4963;
input x_4964;
input x_4965;
input x_4966;
input x_4967;
input x_4968;
input x_4969;
input x_4970;
input x_4971;
input x_4972;
input x_4973;
input x_4974;
input x_4975;
input x_4976;
input x_4977;
input x_4978;
input x_4979;
input x_4980;
input x_4981;
input x_4982;
input x_4983;
input x_4984;
input x_4985;
input x_4986;
input x_4987;
input x_4988;
input x_4989;
input x_4990;
input x_4991;
input x_4992;
input x_4993;
input x_4994;
input x_4995;
input x_4996;
input x_4997;
input x_4998;
input x_4999;
input x_5000;
input x_5001;
input x_5002;
input x_5003;
input x_5004;
input x_5005;
input x_5006;
input x_5007;
input x_5008;
input x_5009;
input x_5010;
input x_5011;
input x_5012;
input x_5013;
input x_5014;
input x_5015;
input x_5016;
input x_5017;
input x_5018;
input x_5019;
input x_5020;
input x_5021;
input x_5022;
input x_5023;
input x_5024;
input x_5025;
input x_5026;
input x_5027;
input x_5028;
input x_5029;
input x_5030;
input x_5031;
input x_5032;
input x_5033;
input x_5034;
input x_5035;
input x_5036;
input x_5037;
input x_5038;
input x_5039;
input x_5040;
input x_5041;
input x_5042;
input x_5043;
input x_5044;
input x_5045;
input x_5046;
input x_5047;
input x_5048;
input x_5049;
input x_5050;
input x_5051;
input x_5052;
input x_5053;
input x_5054;
input x_5055;
input x_5056;
input x_5057;
input x_5058;
input x_5059;
input x_5060;
input x_5061;
input x_5062;
input x_5063;
input x_5064;
input x_5065;
input x_5066;
input x_5067;
input x_5068;
input x_5069;
input x_5070;
input x_5071;
input x_5072;
input x_5073;
input x_5074;
input x_5075;
input x_5076;
input x_5077;
input x_5078;
input x_5079;
input x_5080;
input x_5081;
input x_5082;
input x_5083;
input x_5084;
input x_5085;
input x_5086;
input x_5087;
input x_5088;
input x_5089;
input x_5090;
input x_5091;
input x_5092;
input x_5093;
input x_5094;
input x_5095;
input x_5096;
input x_5097;
input x_5098;
input x_5099;
input x_5100;
input x_5101;
input x_5102;
input x_5103;
input x_5104;
input x_5105;
input x_5106;
input x_5107;
input x_5108;
input x_5109;
input x_5110;
input x_5111;
input x_5112;
input x_5113;
input x_5114;
input x_5115;
input x_5116;
input x_5117;
input x_5118;
input x_5119;
input x_5120;
input x_5121;
input x_5122;
input x_5123;
input x_5124;
input x_5125;
input x_5126;
input x_5127;
input x_5128;
input x_5129;
input x_5130;
input x_5131;
input x_5132;
input x_5133;
input x_5134;
input x_5135;
input x_5136;
input x_5137;
input x_5138;
input x_5139;
input x_5140;
input x_5141;
input x_5142;
input x_5143;
input x_5144;
input x_5145;
input x_5146;
input x_5147;
input x_5148;
input x_5149;
input x_5150;
input x_5151;
input x_5152;
input x_5153;
input x_5154;
input x_5155;
input x_5156;
input x_5157;
input x_5158;
input x_5159;
input x_5160;
input x_5161;
input x_5162;
input x_5163;
input x_5164;
input x_5165;
input x_5166;
input x_5167;
input x_5168;
input x_5169;
input x_5170;
input x_5171;
input x_5172;
input x_5173;
input x_5174;
input x_5175;
input x_5176;
input x_5177;
input x_5178;
input x_5179;
input x_5180;
input x_5181;
input x_5182;
input x_5183;
input x_5184;
input x_5185;
input x_5186;
input x_5187;
input x_5188;
input x_5189;
input x_5190;
input x_5191;
input x_5192;
input x_5193;
input x_5194;
input x_5195;
input x_5196;
input x_5197;
input x_5198;
input x_5199;
input x_5200;
input x_5201;
input x_5202;
input x_5203;
input x_5204;
input x_5205;
input x_5206;
input x_5207;
input x_5208;
input x_5209;
input x_5210;
input x_5211;
input x_5212;
input x_5213;
input x_5214;
input x_5215;
input x_5216;
input x_5217;
input x_5218;
input x_5219;
input x_5220;
input x_5221;
input x_5222;
input x_5223;
input x_5224;
input x_5225;
input x_5226;
input x_5227;
input x_5228;
input x_5229;
input x_5230;
input x_5231;
input x_5232;
input x_5233;
input x_5234;
input x_5235;
input x_5236;
input x_5237;
input x_5238;
input x_5239;
input x_5240;
input x_5241;
input x_5242;
input x_5243;
input x_5244;
input x_5245;
input x_5246;
input x_5247;
input x_5248;
input x_5249;
input x_5250;
input x_5251;
input x_5252;
input x_5253;
input x_5254;
input x_5255;
input x_5256;
input x_5257;
input x_5258;
input x_5259;
input x_5260;
input x_5261;
input x_5262;
input x_5263;
input x_5264;
input x_5265;
input x_5266;
input x_5267;
input x_5268;
input x_5269;
input x_5270;
input x_5271;
input x_5272;
input x_5273;
input x_5274;
input x_5275;
input x_5276;
input x_5277;
input x_5278;
input x_5279;
input x_5280;
input x_5281;
input x_5282;
input x_5283;
input x_5284;
input x_5285;
input x_5286;
input x_5287;
input x_5288;
input x_5289;
input x_5290;
input x_5291;
input x_5292;
input x_5293;
input x_5294;
input x_5295;
input x_5296;
input x_5297;
input x_5298;
input x_5299;
input x_5300;
input x_5301;
input x_5302;
input x_5303;
input x_5304;
input x_5305;
input x_5306;
input x_5307;
input x_5308;
input x_5309;
input x_5310;
input x_5311;
input x_5312;
input x_5313;
input x_5314;
input x_5315;
input x_5316;
input x_5317;
input x_5318;
input x_5319;
input x_5320;
input x_5321;
input x_5322;
input x_5323;
input x_5324;
input x_5325;
input x_5326;
input x_5327;
input x_5328;
input x_5329;
input x_5330;
input x_5331;
input x_5332;
input x_5333;
input x_5334;
input x_5335;
input x_5336;
input x_5337;
input x_5338;
input x_5339;
input x_5340;
input x_5341;
input x_5342;
input x_5343;
input x_5344;
input x_5345;
input x_5346;
input x_5347;
input x_5348;
input x_5349;
input x_5350;
input x_5351;
input x_5352;
input x_5353;
input x_5354;
input x_5355;
input x_5356;
input x_5357;
input x_5358;
input x_5359;
input x_5360;
input x_5361;
input x_5362;
input x_5363;
input x_5364;
input x_5365;
input x_5366;
input x_5367;
input x_5368;
input x_5369;
input x_5370;
input x_5371;
input x_5372;
input x_5373;
input x_5374;
input x_5375;
input x_5376;
input x_5377;
input x_5378;
input x_5379;
input x_5380;
input x_5381;
input x_5382;
input x_5383;
input x_5384;
input x_5385;
input x_5386;
input x_5387;
input x_5388;
input x_5389;
input x_5390;
input x_5391;
input x_5392;
input x_5393;
input x_5394;
input x_5395;
input x_5396;
input x_5397;
input x_5398;
input x_5399;
input x_5400;
input x_5401;
input x_5402;
input x_5403;
input x_5404;
input x_5405;
input x_5406;
input x_5407;
input x_5408;
input x_5409;
input x_5410;
input x_5411;
input x_5412;
input x_5413;
input x_5414;
input x_5415;
input x_5416;
input x_5417;
input x_5418;
input x_5419;
input x_5420;
input x_5421;
input x_5422;
input x_5423;
input x_5424;
input x_5425;
input x_5426;
input x_5427;
input x_5428;
input x_5429;
input x_5430;
input x_5431;
input x_5432;
input x_5433;
input x_5434;
input x_5435;
input x_5436;
input x_5437;
input x_5438;
input x_5439;
input x_5440;
input x_5441;
input x_5442;
input x_5443;
input x_5444;
input x_5445;
input x_5446;
input x_5447;
input x_5448;
input x_5449;
input x_5450;
input x_5451;
input x_5452;
input x_5453;
input x_5454;
input x_5455;
input x_5456;
input x_5457;
input x_5458;
input x_5459;
input x_5460;
input x_5461;
input x_5462;
input x_5463;
input x_5464;
input x_5465;
input x_5466;
input x_5467;
input x_5468;
input x_5469;
input x_5470;
input x_5471;
input x_5472;
input x_5473;
input x_5474;
input x_5475;
input x_5476;
input x_5477;
input x_5478;
input x_5479;
input x_5480;
input x_5481;
input x_5482;
input x_5483;
input x_5484;
input x_5485;
input x_5486;
input x_5487;
input x_5488;
input x_5489;
input x_5490;
input x_5491;
input x_5492;
input x_5493;
input x_5494;
input x_5495;
input x_5496;
input x_5497;
input x_5498;
input x_5499;
input x_5500;
input x_5501;
input x_5502;
input x_5503;
input x_5504;
input x_5505;
input x_5506;
input x_5507;
input x_5508;
input x_5509;
input x_5510;
input x_5511;
input x_5512;
input x_5513;
input x_5514;
input x_5515;
input x_5516;
input x_5517;
input x_5518;
input x_5519;
input x_5520;
input x_5521;
input x_5522;
input x_5523;
input x_5524;
input x_5525;
input x_5526;
input x_5527;
input x_5528;
input x_5529;
input x_5530;
input x_5531;
input x_5532;
input x_5533;
input x_5534;
input x_5535;
input x_5536;
input x_5537;
input x_5538;
input x_5539;
input x_5540;
input x_5541;
input x_5542;
input x_5543;
input x_5544;
input x_5545;
input x_5546;
input x_5547;
input x_5548;
input x_5549;
input x_5550;
input x_5551;
input x_5552;
input x_5553;
input x_5554;
input x_5555;
input x_5556;
input x_5557;
input x_5558;
input x_5559;
input x_5560;
input x_5561;
input x_5562;
input x_5563;
input x_5564;
input x_5565;
input x_5566;
input x_5567;
input x_5568;
input x_5569;
input x_5570;
input x_5571;
input x_5572;
input x_5573;
input x_5574;
input x_5575;
input x_5576;
input x_5577;
input x_5578;
input x_5579;
input x_5580;
input x_5581;
input x_5582;
input x_5583;
input x_5584;
input x_5585;
input x_5586;
input x_5587;
input x_5588;
input x_5589;
input x_5590;
input x_5591;
input x_5592;
input x_5593;
input x_5594;
input x_5595;
input x_5596;
input x_5597;
input x_5598;
input x_5599;
input x_5600;
input x_5601;
input x_5602;
input x_5603;
input x_5604;
input x_5605;
input x_5606;
input x_5607;
input x_5608;
input x_5609;
input x_5610;
input x_5611;
input x_5612;
input x_5613;
input x_5614;
input x_5615;
input x_5616;
input x_5617;
input x_5618;
input x_5619;
input x_5620;
input x_5621;
input x_5622;
input x_5623;
input x_5624;
input x_5625;
input x_5626;
input x_5627;
input x_5628;
input x_5629;
input x_5630;
input x_5631;
input x_5632;
input x_5633;
input x_5634;
input x_5635;
input x_5636;
input x_5637;
input x_5638;
input x_5639;
input x_5640;
input x_5641;
input x_5642;
input x_5643;
input x_5644;
input x_5645;
input x_5646;
input x_5647;
input x_5648;
input x_5649;
input x_5650;
input x_5651;
input x_5652;
input x_5653;
input x_5654;
input x_5655;
input x_5656;
input x_5657;
input x_5658;
input x_5659;
input x_5660;
input x_5661;
input x_5662;
input x_5663;
input x_5664;
input x_5665;
input x_5666;
input x_5667;
input x_5668;
input x_5669;
input x_5670;
input x_5671;
input x_5672;
input x_5673;
input x_5674;
input x_5675;
input x_5676;
input x_5677;
input x_5678;
input x_5679;
input x_5680;
input x_5681;
input x_5682;
input x_5683;
input x_5684;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_2770;
wire n_2771;
wire n_2772;
wire n_2773;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_2790;
wire n_2791;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2796;
wire n_2797;
wire n_2798;
wire n_2799;
wire n_2800;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2808;
wire n_2809;
wire n_2810;
wire n_2811;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2816;
wire n_2817;
wire n_2818;
wire n_2819;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2827;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2832;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2837;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2845;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_2850;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2875;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_2879;
wire n_2880;
wire n_2881;
wire n_2882;
wire n_2883;
wire n_2884;
wire n_2885;
wire n_2886;
wire n_2887;
wire n_2888;
wire n_2889;
wire n_2890;
wire n_2891;
wire n_2892;
wire n_2893;
wire n_2894;
wire n_2895;
wire n_2896;
wire n_2897;
wire n_2898;
wire n_2899;
wire n_2900;
wire n_2901;
wire n_2902;
wire n_2903;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2908;
wire n_2909;
wire n_2910;
wire n_2911;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2923;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2928;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2944;
wire n_2945;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_3069;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_3400;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_3410;
wire n_3411;
wire n_3412;
wire n_3413;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_3428;
wire n_3429;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4038;
wire n_4039;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4125;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire n_4159;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_4178;
wire n_4179;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_4187;
wire n_4188;
wire n_4189;
wire n_4190;
wire n_4191;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_4200;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4216;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_4240;
wire n_4241;
wire n_4242;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire n_4285;
wire n_4286;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4348;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_4790;
wire n_4791;
wire n_4792;
wire n_4793;
wire n_4794;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4803;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4854;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4865;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4876;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4882;
wire n_4883;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire n_4888;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4893;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4898;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4910;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4924;
wire n_4925;
wire n_4926;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_4930;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4934;
wire n_4935;
wire n_4936;
wire n_4937;
wire n_4938;
wire n_4939;
wire n_4940;
wire n_4941;
wire n_4942;
wire n_4943;
wire n_4944;
wire n_4945;
wire n_4946;
wire n_4947;
wire n_4948;
wire n_4949;
wire n_4950;
wire n_4951;
wire n_4952;
wire n_4953;
wire n_4954;
wire n_4955;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_4960;
wire n_4961;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4967;
wire n_4968;
wire n_4969;
wire n_4970;
wire n_4971;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4977;
wire n_4978;
wire n_4979;
wire n_4980;
wire n_4981;
wire n_4982;
wire n_4983;
wire n_4984;
wire n_4985;
wire n_4986;
wire n_4987;
wire n_4988;
wire n_4989;
wire n_4990;
wire n_4991;
wire n_4992;
wire n_4993;
wire n_4994;
wire n_4995;
wire n_4996;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_5000;
wire n_5001;
wire n_5002;
wire n_5003;
wire n_5004;
wire n_5005;
wire n_5006;
wire n_5007;
wire n_5008;
wire n_5009;
wire n_5010;
wire n_5011;
wire n_5012;
wire n_5013;
wire n_5014;
wire n_5015;
wire n_5016;
wire n_5017;
wire n_5018;
wire n_5019;
wire n_5020;
wire n_5021;
wire n_5022;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5027;
wire n_5028;
wire n_5029;
wire n_5030;
wire n_5031;
wire n_5032;
wire n_5033;
wire n_5034;
wire n_5035;
wire n_5036;
wire n_5037;
wire n_5038;
wire n_5039;
wire n_5040;
wire n_5041;
wire n_5042;
wire n_5043;
wire n_5044;
wire n_5045;
wire n_5046;
wire n_5047;
wire n_5048;
wire n_5049;
wire n_5050;
wire n_5051;
wire n_5052;
wire n_5053;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_5058;
wire n_5059;
wire n_5060;
wire n_5061;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5066;
wire n_5067;
wire n_5068;
wire n_5069;
wire n_5070;
wire n_5071;
wire n_5072;
wire n_5073;
wire n_5074;
wire n_5075;
wire n_5076;
wire n_5077;
wire n_5078;
wire n_5079;
wire n_5080;
wire n_5081;
wire n_5082;
wire n_5083;
wire n_5084;
wire n_5085;
wire n_5086;
wire n_5087;
wire n_5088;
wire n_5089;
wire n_5090;
wire n_5091;
wire n_5092;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire n_5097;
wire n_5098;
wire n_5099;
wire n_5100;
wire n_5101;
wire n_5102;
wire n_5103;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5118;
wire n_5119;
wire n_5120;
wire n_5121;
wire n_5122;
wire n_5123;
wire n_5124;
wire n_5125;
wire n_5126;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5133;
wire n_5134;
wire n_5135;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire n_5148;
wire n_5149;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5155;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_5160;
wire n_5161;
wire n_5162;
wire n_5163;
wire n_5164;
wire n_5165;
wire n_5166;
wire n_5167;
wire n_5168;
wire n_5169;
wire n_5170;
wire n_5171;
wire n_5172;
wire n_5173;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_5179;
wire n_5180;
wire n_5181;
wire n_5182;
wire n_5183;
wire n_5184;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_5190;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_5200;
wire n_5201;
wire n_5202;
wire n_5203;
wire n_5204;
wire n_5205;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5214;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_5219;
wire n_5220;
wire n_5221;
wire n_5222;
wire n_5223;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_5237;
wire n_5238;
wire n_5239;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5245;
wire n_5246;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_5250;
wire n_5251;
wire n_5252;
wire n_5253;
wire n_5254;
wire n_5255;
wire n_5256;
wire n_5257;
wire n_5258;
wire n_5259;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5264;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_5268;
wire n_5269;
wire n_5270;
wire n_5271;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5278;
wire n_5279;
wire n_5280;
wire n_5281;
wire n_5282;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_5290;
wire n_5291;
wire n_5292;
wire n_5293;
wire n_5294;
wire n_5295;
wire n_5296;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_5300;
wire n_5301;
wire n_5302;
wire n_5303;
wire n_5304;
wire n_5305;
wire n_5306;
wire n_5307;
wire n_5308;
wire n_5309;
wire n_5310;
wire n_5311;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire n_5317;
wire n_5318;
wire n_5319;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5326;
wire n_5327;
wire n_5328;
wire n_5329;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5337;
wire n_5338;
wire n_5339;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5347;
wire n_5348;
wire n_5349;
wire n_5350;
wire n_5351;
wire n_5352;
wire n_5353;
wire n_5354;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_5360;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5366;
wire n_5367;
wire n_5368;
wire n_5369;
wire n_5370;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5376;
wire n_5377;
wire n_5378;
wire n_5379;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5383;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire n_5388;
wire n_5389;
wire n_5390;
wire n_5391;
wire n_5392;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5396;
wire n_5397;
wire n_5398;
wire n_5399;
wire n_5400;
wire n_5401;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire n_5407;
wire n_5408;
wire n_5409;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5413;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_5419;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5427;
wire n_5428;
wire n_5429;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire n_5435;
wire n_5436;
wire n_5437;
wire n_5438;
wire n_5439;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5445;
wire n_5446;
wire n_5447;
wire n_5448;
wire n_5449;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5453;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5466;
wire n_5467;
wire n_5468;
wire n_5469;
wire n_5470;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5474;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_5479;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_5490;
wire n_5491;
wire n_5492;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5507;
wire n_5508;
wire n_5509;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5513;
wire n_5514;
wire n_5515;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5519;
wire n_5520;
wire n_5521;
wire n_5522;
wire n_5523;
wire n_5524;
wire n_5525;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5533;
wire n_5534;
wire n_5535;
wire n_5536;
wire n_5537;
wire n_5538;
wire n_5539;
wire n_5540;
wire n_5541;
wire n_5542;
wire n_5543;
wire n_5544;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5560;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5585;
wire n_5586;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_5590;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5597;
wire n_5598;
wire n_5599;
wire n_5600;
wire n_5601;
wire n_5602;
wire n_5603;
wire n_5604;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5615;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5623;
wire n_5624;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire n_5645;
wire n_5646;
wire n_5647;
wire n_5648;
wire n_5649;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5653;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire n_5668;
wire n_5669;
wire n_5670;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5678;
wire n_5679;
wire n_5680;
wire n_5681;
wire n_5682;
wire n_5683;
wire n_5684;
wire n_5685;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5694;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_5699;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5711;
wire n_5712;
wire n_5713;
wire n_5714;
wire n_5715;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_5720;
wire n_5721;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5729;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5734;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5738;
wire n_5739;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5746;
wire n_5747;
wire n_5748;
wire n_5749;
wire n_5750;
wire n_5751;
wire n_5752;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5758;
wire n_5759;
wire n_5760;
wire n_5761;
wire n_5762;
wire n_5763;
wire n_5764;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5771;
wire n_5772;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_5780;
wire n_5781;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_5790;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5794;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire n_5799;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5803;
wire n_5804;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_5809;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5817;
wire n_5818;
wire n_5819;
wire n_5820;
wire n_5821;
wire n_5822;
wire n_5823;
wire n_5824;
wire n_5825;
wire n_5826;
wire n_5827;
wire n_5828;
wire n_5829;
wire n_5830;
wire n_5831;
wire n_5832;
wire n_5833;
wire n_5834;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5843;
wire n_5844;
wire n_5845;
wire n_5846;
wire n_5847;
wire n_5848;
wire n_5849;
wire n_5850;
wire n_5851;
wire n_5852;
wire n_5853;
wire n_5854;
wire n_5855;
wire n_5856;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5865;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_5869;
wire n_5870;
wire n_5871;
wire n_5872;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire n_5885;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_5890;
wire n_5891;
wire n_5892;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5903;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5908;
wire n_5909;
wire n_5910;
wire n_5911;
wire n_5912;
wire n_5913;
wire n_5914;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire n_5920;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_5930;
wire n_5931;
wire n_5932;
wire n_5933;
wire n_5934;
wire n_5935;
wire n_5936;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_5940;
wire n_5941;
wire n_5942;
wire n_5943;
wire n_5944;
wire n_5945;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5954;
wire n_5955;
wire n_5956;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_5960;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_5970;
wire n_5971;
wire n_5972;
wire n_5973;
wire n_5974;
wire n_5975;
wire n_5976;
wire n_5977;
wire n_5978;
wire n_5979;
wire n_5980;
wire n_5981;
wire n_5982;
wire n_5983;
wire n_5984;
wire n_5985;
wire n_5986;
wire n_5987;
wire n_5988;
wire n_5989;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5993;
wire n_5994;
wire n_5995;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_6000;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire n_6014;
wire n_6015;
wire n_6016;
wire n_6017;
wire n_6018;
wire n_6019;
wire n_6020;
wire n_6021;
wire n_6022;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6027;
wire n_6028;
wire n_6029;
wire n_6030;
wire n_6031;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6035;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_6039;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6045;
wire n_6046;
wire n_6047;
wire n_6048;
wire n_6049;
wire n_6050;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire n_6056;
wire n_6057;
wire n_6058;
wire n_6059;
wire n_6060;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_6070;
wire n_6071;
wire n_6072;
wire n_6073;
wire n_6074;
wire n_6075;
wire n_6076;
wire n_6077;
wire n_6078;
wire n_6079;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire n_6084;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6088;
wire n_6089;
wire n_6090;
wire n_6091;
wire n_6092;
wire n_6093;
wire n_6094;
wire n_6095;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_6099;
wire n_6100;
wire n_6101;
wire n_6102;
wire n_6103;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_6110;
wire n_6111;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_6120;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6126;
wire n_6127;
wire n_6128;
wire n_6129;
wire n_6130;
wire n_6131;
wire n_6132;
wire n_6133;
wire n_6134;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_6150;
wire n_6151;
wire n_6152;
wire n_6153;
wire n_6154;
wire n_6155;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_6160;
wire n_6161;
wire n_6162;
wire n_6163;
wire n_6164;
wire n_6165;
wire n_6166;
wire n_6167;
wire n_6168;
wire n_6169;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6174;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_6190;
wire n_6191;
wire n_6192;
wire n_6193;
wire n_6194;
wire n_6195;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_6199;
wire n_6200;
wire n_6201;
wire n_6202;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_6210;
wire n_6211;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6216;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_6220;
wire n_6221;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6227;
wire n_6228;
wire n_6229;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6236;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_6240;
wire n_6241;
wire n_6242;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6246;
wire n_6247;
wire n_6248;
wire n_6249;
wire n_6250;
wire n_6251;
wire n_6252;
wire n_6253;
wire n_6254;
wire n_6255;
wire n_6256;
wire n_6257;
wire n_6258;
wire n_6259;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6264;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_6270;
wire n_6271;
wire n_6272;
wire n_6273;
wire n_6274;
wire n_6275;
wire n_6276;
wire n_6277;
wire n_6278;
wire n_6279;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6283;
wire n_6284;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_6289;
wire n_6290;
wire n_6291;
wire n_6292;
wire n_6293;
wire n_6294;
wire n_6295;
wire n_6296;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_6300;
wire n_6301;
wire n_6302;
wire n_6303;
wire n_6304;
wire n_6305;
wire n_6306;
wire n_6307;
wire n_6308;
wire n_6309;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6314;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_6320;
wire n_6321;
wire n_6322;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_6330;
wire n_6331;
wire n_6332;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6336;
wire n_6337;
wire n_6338;
wire n_6339;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire n_6344;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire n_6349;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_6360;
wire n_6361;
wire n_6362;
wire n_6363;
wire n_6364;
wire n_6365;
wire n_6366;
wire n_6367;
wire n_6368;
wire n_6369;
wire n_6370;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6375;
wire n_6376;
wire n_6377;
wire n_6378;
wire n_6379;
wire n_6380;
wire n_6381;
wire n_6382;
wire n_6383;
wire n_6384;
wire n_6385;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire n_6397;
wire n_6398;
wire n_6399;
wire n_6400;
wire n_6401;
wire n_6402;
wire n_6403;
wire n_6404;
wire n_6405;
wire n_6406;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_6410;
wire n_6411;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire n_6417;
wire n_6418;
wire n_6419;
wire n_6420;
wire n_6421;
wire n_6422;
wire n_6423;
wire n_6424;
wire n_6425;
wire n_6426;
wire n_6427;
wire n_6428;
wire n_6429;
wire n_6430;
wire n_6431;
wire n_6432;
wire n_6433;
wire n_6434;
wire n_6435;
wire n_6436;
wire n_6437;
wire n_6438;
wire n_6439;
wire n_6440;
wire n_6441;
wire n_6442;
wire n_6443;
wire n_6444;
wire n_6445;
wire n_6446;
wire n_6447;
wire n_6448;
wire n_6449;
wire n_6450;
wire n_6451;
wire n_6452;
wire n_6453;
wire n_6454;
wire n_6455;
wire n_6456;
wire n_6457;
wire n_6458;
wire n_6459;
wire n_6460;
wire n_6461;
wire n_6462;
wire n_6463;
wire n_6464;
wire n_6465;
wire n_6466;
wire n_6467;
wire n_6468;
wire n_6469;
wire n_6470;
wire n_6471;
wire n_6472;
wire n_6473;
wire n_6474;
wire n_6475;
wire n_6476;
wire n_6477;
wire n_6478;
wire n_6479;
wire n_6480;
wire n_6481;
wire n_6482;
wire n_6483;
wire n_6484;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_6490;
wire n_6491;
wire n_6492;
wire n_6493;
wire n_6494;
wire n_6495;
wire n_6496;
wire n_6497;
wire n_6498;
wire n_6499;
wire n_6500;
wire n_6501;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6508;
wire n_6509;
wire n_6510;
wire n_6511;
wire n_6512;
wire n_6513;
wire n_6514;
wire n_6515;
wire n_6516;
wire n_6517;
wire n_6518;
wire n_6519;
wire n_6520;
wire n_6521;
wire n_6522;
wire n_6523;
wire n_6524;
wire n_6525;
wire n_6526;
wire n_6527;
wire n_6528;
wire n_6529;
wire n_6530;
wire n_6531;
wire n_6532;
wire n_6533;
wire n_6534;
wire n_6535;
wire n_6536;
wire n_6537;
wire n_6538;
wire n_6539;
wire n_6540;
wire n_6541;
wire n_6542;
wire n_6543;
wire n_6544;
wire n_6545;
wire n_6546;
wire n_6547;
wire n_6548;
wire n_6549;
wire n_6550;
wire n_6551;
wire n_6552;
wire n_6553;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_6559;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6566;
wire n_6567;
wire n_6568;
wire n_6569;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6573;
wire n_6574;
wire n_6575;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6584;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6588;
wire n_6589;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_6600;
wire n_6601;
wire n_6602;
wire n_6603;
wire n_6604;
wire n_6605;
wire n_6606;
wire n_6607;
wire n_6608;
wire n_6609;
wire n_6610;
wire n_6611;
wire n_6612;
wire n_6613;
wire n_6614;
wire n_6615;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_6620;
wire n_6621;
wire n_6622;
wire n_6623;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_6629;
wire n_6630;
wire n_6631;
wire n_6632;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6636;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6647;
wire n_6648;
wire n_6649;
wire n_6650;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6657;
wire n_6658;
wire n_6659;
wire n_6660;
wire n_6661;
wire n_6662;
wire n_6663;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6677;
wire n_6678;
wire n_6679;
wire n_6680;
wire n_6681;
wire n_6682;
wire n_6683;
wire n_6684;
wire n_6685;
wire n_6686;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_6690;
wire n_6691;
wire n_6692;
wire n_6693;
wire n_6694;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_6699;
wire n_6700;
wire n_6701;
wire n_6702;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_6709;
wire n_6710;
wire n_6711;
wire n_6712;
wire n_6713;
wire n_6714;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6726;
wire n_6727;
wire n_6728;
wire n_6729;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6735;
wire n_6736;
wire n_6737;
wire n_6738;
wire n_6739;
wire n_6740;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6744;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_6750;
wire n_6751;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6757;
wire n_6758;
wire n_6759;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6766;
wire n_6767;
wire n_6768;
wire n_6769;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire n_6777;
wire n_6778;
wire n_6779;
wire n_6780;
wire n_6781;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6785;
wire n_6786;
wire n_6787;
wire n_6788;
wire n_6789;
wire n_6790;
wire n_6791;
wire n_6792;
wire n_6793;
wire n_6794;
wire n_6795;
wire n_6796;
wire n_6797;
wire n_6798;
wire n_6799;
wire n_6800;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6805;
wire n_6806;
wire n_6807;
wire n_6808;
wire n_6809;
wire n_6810;
wire n_6811;
wire n_6812;
wire n_6813;
wire n_6814;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_6820;
wire n_6821;
wire n_6822;
wire n_6823;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6827;
wire n_6828;
wire n_6829;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_6837;
wire n_6838;
wire n_6839;
wire n_6840;
wire n_6841;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6846;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6888;
wire n_6889;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6894;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_6900;
wire n_6901;
wire n_6902;
wire n_6903;
wire n_6904;
wire n_6905;
wire n_6906;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_6910;
wire n_6911;
wire n_6912;
wire n_6913;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6917;
wire n_6918;
wire n_6919;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_6930;
wire n_6931;
wire n_6932;
wire n_6933;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6954;
wire n_6955;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_6970;
wire n_6971;
wire n_6972;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6978;
wire n_6979;
wire n_6980;
wire n_6981;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7018;
wire n_7019;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire n_7076;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7104;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7115;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire n_7125;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_7130;
wire n_7131;
wire n_7132;
wire n_7133;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_7140;
wire n_7141;
wire n_7142;
wire n_7143;
wire n_7144;
wire n_7145;
wire n_7146;
wire n_7147;
wire n_7148;
wire n_7149;
wire n_7150;
wire n_7151;
wire n_7152;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7174;
wire n_7175;
wire n_7176;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_7180;
wire n_7181;
wire n_7182;
wire n_7183;
wire n_7184;
wire n_7185;
wire n_7186;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_7190;
wire n_7191;
wire n_7192;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_7200;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7205;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_7220;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7230;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_7319;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7325;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7336;
wire n_7337;
wire n_7338;
wire n_7339;
wire n_7340;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_7350;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7367;
wire n_7368;
wire n_7369;
wire n_7370;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_7380;
wire n_7381;
wire n_7382;
wire n_7383;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_7390;
wire n_7391;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7504;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7533;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7553;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7641;
wire n_7642;
wire n_7643;
wire n_7644;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7688;
wire n_7689;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7694;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire n_7729;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7758;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7770;
wire n_7771;
wire n_7772;
wire n_7773;
wire n_7774;
wire n_7775;
wire n_7776;
wire n_7777;
wire n_7778;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7825;
wire n_7826;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7833;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7837;
wire n_7838;
wire n_7839;
wire n_7840;
wire n_7841;
wire n_7842;
wire n_7843;
wire n_7844;
wire n_7845;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire n_7850;
wire n_7851;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7856;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7867;
wire n_7868;
wire n_7869;
wire n_7870;
wire n_7871;
wire n_7872;
wire n_7873;
wire n_7874;
wire n_7875;
wire n_7876;
wire n_7877;
wire n_7878;
wire n_7879;
wire n_7880;
wire n_7881;
wire n_7882;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7886;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_7890;
wire n_7891;
wire n_7892;
wire n_7893;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_7899;
wire n_7900;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_7904;
wire n_7905;
wire n_7906;
wire n_7907;
wire n_7908;
wire n_7909;
wire n_7910;
wire n_7911;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire n_7926;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_7930;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_7940;
wire n_7941;
wire n_7942;
wire n_7943;
wire n_7944;
wire n_7945;
wire n_7946;
wire n_7947;
wire n_7948;
wire n_7949;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7956;
wire n_7957;
wire n_7958;
wire n_7959;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_7970;
wire n_7971;
wire n_7972;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_7980;
wire n_7981;
wire n_7982;
wire n_7983;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7994;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_8000;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8013;
wire n_8014;
wire n_8015;
wire n_8016;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_8020;
wire n_8021;
wire n_8022;
wire n_8023;
wire n_8024;
wire n_8025;
wire n_8026;
wire n_8027;
wire n_8028;
wire n_8029;
wire n_8030;
wire n_8031;
wire n_8032;
wire n_8033;
wire n_8034;
wire n_8035;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_8049;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8055;
wire n_8056;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_8060;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_8070;
wire n_8071;
wire n_8072;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8076;
wire n_8077;
wire n_8078;
wire n_8079;
wire n_8080;
wire n_8081;
wire n_8082;
wire n_8083;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_8088;
wire n_8089;
wire n_8090;
wire n_8091;
wire n_8092;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_8110;
wire n_8111;
wire n_8112;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8116;
wire n_8117;
wire n_8118;
wire n_8119;
wire n_8120;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_8129;
wire n_8130;
wire n_8131;
wire n_8132;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8137;
wire n_8138;
wire n_8139;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire n_8146;
wire n_8147;
wire n_8148;
wire n_8149;
wire n_8150;
wire n_8151;
wire n_8152;
wire n_8153;
wire n_8154;
wire n_8155;
wire n_8156;
wire n_8157;
wire n_8158;
wire n_8159;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire n_8164;
wire n_8165;
wire n_8166;
wire n_8167;
wire n_8168;
wire n_8169;
wire n_8170;
wire n_8171;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire n_8178;
wire n_8179;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire n_8184;
wire n_8185;
wire n_8186;
wire n_8187;
wire n_8188;
wire n_8189;
wire n_8190;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8194;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8198;
wire n_8199;
wire n_8200;
wire n_8201;
wire n_8202;
wire n_8203;
wire n_8204;
wire n_8205;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_8209;
wire n_8210;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8214;
wire n_8215;
wire n_8216;
wire n_8217;
wire n_8218;
wire n_8219;
wire n_8220;
wire n_8221;
wire n_8222;
wire n_8223;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8228;
wire n_8229;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8233;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_8240;
wire n_8241;
wire n_8242;
wire n_8243;
wire n_8244;
wire n_8245;
wire n_8246;
wire n_8247;
wire n_8248;
wire n_8249;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8253;
wire n_8254;
wire n_8255;
wire n_8256;
wire n_8257;
wire n_8258;
wire n_8259;
wire n_8260;
wire n_8261;
wire n_8262;
wire n_8263;
wire n_8264;
wire n_8265;
wire n_8266;
wire n_8267;
wire n_8268;
wire n_8269;
wire n_8270;
wire n_8271;
wire n_8272;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8276;
wire n_8277;
wire n_8278;
wire n_8279;
wire n_8280;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8286;
wire n_8287;
wire n_8288;
wire n_8289;
wire n_8290;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire n_8297;
wire n_8298;
wire n_8299;
wire n_8300;
wire n_8301;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8308;
wire n_8309;
wire n_8310;
wire n_8311;
wire n_8312;
wire n_8313;
wire n_8314;
wire n_8315;
wire n_8316;
wire n_8317;
wire n_8318;
wire n_8319;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8323;
wire n_8324;
wire n_8325;
wire n_8326;
wire n_8327;
wire n_8328;
wire n_8329;
wire n_8330;
wire n_8331;
wire n_8332;
wire n_8333;
wire n_8334;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_8338;
wire n_8339;
wire n_8340;
wire n_8341;
wire n_8342;
wire n_8343;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8347;
wire n_8348;
wire n_8349;
wire n_8350;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8356;
wire n_8357;
wire n_8358;
wire n_8359;
wire n_8360;
wire n_8361;
wire n_8362;
wire n_8363;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8377;
wire n_8378;
wire n_8379;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8383;
wire n_8384;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_8390;
wire n_8391;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8397;
wire n_8398;
wire n_8399;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8408;
wire n_8409;
wire n_8410;
wire n_8411;
wire n_8412;
wire n_8413;
wire n_8414;
wire n_8415;
wire n_8416;
wire n_8417;
wire n_8418;
wire n_8419;
wire n_8420;
wire n_8421;
wire n_8422;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_8470;
wire n_8471;
wire n_8472;
wire n_8473;
wire n_8474;
wire n_8475;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_8500;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8537;
wire n_8538;
wire n_8539;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8543;
wire n_8544;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8577;
wire n_8578;
wire n_8579;
wire n_8580;
wire n_8581;
wire n_8582;
wire n_8583;
wire n_8584;
wire n_8585;
wire n_8586;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8592;
wire n_8593;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8599;
wire n_8600;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_8610;
wire n_8611;
wire n_8612;
wire n_8613;
wire n_8614;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8654;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8663;
wire n_8664;
wire n_8665;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_8669;
wire n_8670;
wire n_8671;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_8679;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8683;
wire n_8684;
wire n_8685;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_8690;
wire n_8691;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8696;
wire n_8697;
wire n_8698;
wire n_8699;
wire n_8700;
wire n_8701;
wire n_8702;
wire n_8703;
wire n_8704;
wire n_8705;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_8710;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8715;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_8720;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8738;
wire n_8739;
wire n_8740;
wire n_8741;
wire n_8742;
wire n_8743;
wire n_8744;
wire n_8745;
wire n_8746;
wire n_8747;
wire n_8748;
wire n_8749;
wire n_8750;
wire n_8751;
wire n_8752;
wire n_8753;
wire n_8754;
wire n_8755;
wire n_8756;
wire n_8757;
wire n_8758;
wire n_8759;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8763;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8768;
wire n_8769;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_8777;
wire n_8778;
wire n_8779;
wire n_8780;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8785;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_8789;
wire n_8790;
wire n_8791;
wire n_8792;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8796;
wire n_8797;
wire n_8798;
wire n_8799;
wire n_8800;
wire n_8801;
wire n_8802;
wire n_8803;
wire n_8804;
wire n_8805;
wire n_8806;
wire n_8807;
wire n_8808;
wire n_8809;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8814;
wire n_8815;
wire n_8816;
wire n_8817;
wire n_8818;
wire n_8819;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8823;
wire n_8824;
wire n_8825;
wire n_8826;
wire n_8827;
wire n_8828;
wire n_8829;
wire n_8830;
wire n_8831;
wire n_8832;
wire n_8833;
wire n_8834;
wire n_8835;
wire n_8836;
wire n_8837;
wire n_8838;
wire n_8839;
wire n_8840;
wire n_8841;
wire n_8842;
wire n_8843;
wire n_8844;
wire n_8845;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8856;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8866;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_8870;
wire n_8871;
wire n_8872;
wire n_8873;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8878;
wire n_8879;
wire n_8880;
wire n_8881;
wire n_8882;
wire n_8883;
wire n_8884;
wire n_8885;
wire n_8886;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_8890;
wire n_8891;
wire n_8892;
wire n_8893;
wire n_8894;
wire n_8895;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_8900;
wire n_8901;
wire n_8902;
wire n_8903;
wire n_8904;
wire n_8905;
wire n_8906;
wire n_8907;
wire n_8908;
wire n_8909;
wire n_8910;
wire n_8911;
wire n_8912;
wire n_8913;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8917;
wire n_8918;
wire n_8919;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8924;
wire n_8925;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_8929;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8935;
wire n_8936;
wire n_8937;
wire n_8938;
wire n_8939;
wire n_8940;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8948;
wire n_8949;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8956;
wire n_8957;
wire n_8958;
wire n_8959;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_8975;
wire n_8976;
wire n_8977;
wire n_8978;
wire n_8979;
wire n_8980;
wire n_8981;
wire n_8982;
wire n_8983;
wire n_8984;
wire n_8985;
wire n_8986;
wire n_8987;
wire n_8988;
wire n_8989;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_9050;
wire n_9051;
wire n_9052;
wire n_9053;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_9060;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire n_9068;
wire n_9069;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9147;
wire n_9148;
wire n_9149;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_9156;
wire n_9157;
wire n_9158;
wire n_9159;
wire n_9160;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9164;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9186;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_9190;
wire n_9191;
wire n_9192;
wire n_9193;
wire n_9194;
wire n_9195;
wire n_9196;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_9210;
wire n_9211;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9244;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_9248;
wire n_9249;
wire n_9250;
wire n_9251;
wire n_9252;
wire n_9253;
wire n_9254;
wire n_9255;
wire n_9256;
wire n_9257;
wire n_9258;
wire n_9259;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9273;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_9277;
wire n_9278;
wire n_9279;
wire n_9280;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_9288;
wire n_9289;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_9300;
wire n_9301;
wire n_9302;
wire n_9303;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9308;
wire n_9309;
wire n_9310;
wire n_9311;
wire n_9312;
wire n_9313;
wire n_9314;
wire n_9315;
wire n_9316;
wire n_9317;
wire n_9318;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9337;
wire n_9338;
wire n_9339;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_9349;
wire n_9350;
wire n_9351;
wire n_9352;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire n_9358;
wire n_9359;
wire n_9360;
wire n_9361;
wire n_9362;
wire n_9363;
wire n_9364;
wire n_9365;
wire n_9366;
wire n_9367;
wire n_9368;
wire n_9369;
wire n_9370;
wire n_9371;
wire n_9372;
wire n_9373;
wire n_9374;
wire n_9375;
wire n_9376;
wire n_9377;
wire n_9378;
wire n_9379;
wire n_9380;
wire n_9381;
wire n_9382;
wire n_9383;
wire n_9384;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9388;
wire n_9389;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9394;
wire n_9395;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_9410;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9417;
wire n_9418;
wire n_9419;
wire n_9420;
wire n_9421;
wire n_9422;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_9429;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9533;
wire n_9534;
wire n_9535;
wire n_9536;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9566;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9575;
wire n_9576;
wire n_9577;
wire n_9578;
wire n_9579;
wire n_9580;
wire n_9581;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_9589;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9597;
wire n_9598;
wire n_9599;
wire n_9600;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire n_9608;
wire n_9609;
wire n_9610;
wire n_9611;
wire n_9612;
wire n_9613;
wire n_9614;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_9619;
wire n_9620;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_9630;
wire n_9631;
wire n_9632;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9636;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9645;
wire n_9646;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_9650;
wire n_9651;
wire n_9652;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_9660;
wire n_9661;
wire n_9662;
wire n_9663;
wire n_9664;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_9669;
wire n_9670;
wire n_9671;
wire n_9672;
wire n_9673;
wire n_9674;
wire n_9675;
wire n_9676;
wire n_9677;
wire n_9678;
wire n_9679;
wire n_9680;
wire n_9681;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9688;
wire n_9689;
wire n_9690;
wire n_9691;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9695;
wire n_9696;
wire n_9697;
wire n_9698;
wire n_9699;
wire n_9700;
wire n_9701;
wire n_9702;
wire n_9703;
wire n_9704;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9715;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9725;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_9730;
wire n_9731;
wire n_9732;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9736;
wire n_9737;
wire n_9738;
wire n_9739;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9743;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire n_9749;
wire n_9750;
wire n_9751;
wire n_9752;
wire n_9753;
wire n_9754;
wire n_9755;
wire n_9756;
wire n_9757;
wire n_9758;
wire n_9759;
wire n_9760;
wire n_9761;
wire n_9762;
wire n_9763;
wire n_9764;
wire n_9765;
wire n_9766;
wire n_9767;
wire n_9768;
wire n_9769;
wire n_9770;
wire n_9771;
wire n_9772;
wire n_9773;
wire n_9774;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_9778;
wire n_9779;
wire n_9780;
wire n_9781;
wire n_9782;
wire n_9783;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_9790;
wire n_9791;
wire n_9792;
wire n_9793;
wire n_9794;
wire n_9795;
wire n_9796;
wire n_9797;
wire n_9798;
wire n_9799;
wire n_9800;
wire n_9801;
wire n_9802;
wire n_9803;
wire n_9804;
wire n_9805;
wire n_9806;
wire n_9807;
wire n_9808;
wire n_9809;
wire n_9810;
wire n_9811;
wire n_9812;
wire n_9813;
wire n_9814;
wire n_9815;
wire n_9816;
wire n_9817;
wire n_9818;
wire n_9819;
wire n_9820;
wire n_9821;
wire n_9822;
wire n_9823;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9833;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire n_9846;
wire n_9847;
wire n_9848;
wire n_9849;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9863;
wire n_9864;
wire n_9865;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_9870;
wire n_9871;
wire n_9872;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire n_9879;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_9890;
wire n_9891;
wire n_9892;
wire n_9893;
wire n_9894;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_9900;
wire n_9901;
wire n_9902;
wire n_9903;
wire n_9904;
wire n_9905;
wire n_9906;
wire n_9907;
wire n_9908;
wire n_9909;
wire n_9910;
wire n_9911;
wire n_9912;
wire n_9913;
wire n_9914;
wire n_9915;
wire n_9916;
wire n_9917;
wire n_9918;
wire n_9919;
wire n_9920;
wire n_9921;
wire n_9922;
wire n_9923;
wire n_9924;
wire n_9925;
wire n_9926;
wire n_9927;
wire n_9928;
wire n_9929;
wire n_9930;
wire n_9931;
wire n_9932;
wire n_9933;
wire n_9934;
wire n_9935;
wire n_9936;
wire n_9937;
wire n_9938;
wire n_9939;
wire n_9940;
wire n_9941;
wire n_9942;
wire n_9943;
wire n_9944;
wire n_9945;
wire n_9946;
wire n_9947;
wire n_9948;
wire n_9949;
wire n_9950;
wire n_9951;
wire n_9952;
wire n_9953;
wire n_9954;
wire n_9955;
wire n_9956;
wire n_9957;
wire n_9958;
wire n_9959;
wire n_9960;
wire n_9961;
wire n_9962;
wire n_9963;
wire n_9964;
wire n_9965;
wire n_9966;
wire n_9967;
wire n_9968;
wire n_9969;
wire n_9970;
wire n_9971;
wire n_9972;
wire n_9973;
wire n_9974;
wire n_9975;
wire n_9976;
wire n_9977;
wire n_9978;
wire n_9979;
wire n_9980;
wire n_9981;
wire n_9982;
wire n_9983;
wire n_9984;
wire n_9985;
wire n_9986;
wire n_9987;
wire n_9988;
wire n_9989;
wire n_9990;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9994;
wire n_9995;
wire n_9996;
wire n_9997;
wire n_9998;
wire n_9999;
wire n_10000;
wire n_10001;
wire n_10002;
wire n_10003;
wire n_10004;
wire n_10005;
wire n_10006;
wire n_10007;
wire n_10008;
wire n_10009;
wire n_10010;
wire n_10011;
wire n_10012;
wire n_10013;
wire n_10014;
wire n_10015;
wire n_10016;
wire n_10017;
wire n_10018;
wire n_10019;
wire n_10020;
wire n_10021;
wire n_10022;
wire n_10023;
wire n_10024;
wire n_10025;
wire n_10026;
wire n_10027;
wire n_10028;
wire n_10029;
wire n_10030;
wire n_10031;
wire n_10032;
wire n_10033;
wire n_10034;
wire n_10035;
wire n_10036;
wire n_10037;
wire n_10038;
wire n_10039;
wire n_10040;
wire n_10041;
wire n_10042;
wire n_10043;
wire n_10044;
wire n_10045;
wire n_10046;
wire n_10047;
wire n_10048;
wire n_10049;
wire n_10050;
wire n_10051;
wire n_10052;
wire n_10053;
wire n_10054;
wire n_10055;
wire n_10056;
wire n_10057;
wire n_10058;
wire n_10059;
wire n_10060;
wire n_10061;
wire n_10062;
wire n_10063;
wire n_10064;
wire n_10065;
wire n_10066;
wire n_10067;
wire n_10068;
wire n_10069;
wire n_10070;
wire n_10071;
wire n_10072;
wire n_10073;
wire n_10074;
wire n_10075;
wire n_10076;
wire n_10077;
wire n_10078;
wire n_10079;
wire n_10080;
wire n_10081;
wire n_10082;
wire n_10083;
wire n_10084;
wire n_10085;
wire n_10086;
wire n_10087;
wire n_10088;
wire n_10089;
wire n_10090;
wire n_10091;
wire n_10092;
wire n_10093;
wire n_10094;
wire n_10095;
wire n_10096;
wire n_10097;
wire n_10098;
wire n_10099;
wire n_10100;
wire n_10101;
wire n_10102;
wire n_10103;
wire n_10104;
wire n_10105;
wire n_10106;
wire n_10107;
wire n_10108;
wire n_10109;
wire n_10110;
wire n_10111;
wire n_10112;
wire n_10113;
wire n_10114;
wire n_10115;
wire n_10116;
wire n_10117;
wire n_10118;
wire n_10119;
wire n_10120;
wire n_10121;
wire n_10122;
wire n_10123;
wire n_10124;
wire n_10125;
wire n_10126;
wire n_10127;
wire n_10128;
wire n_10129;
wire n_10130;
wire n_10131;
wire n_10132;
wire n_10133;
wire n_10134;
wire n_10135;
wire n_10136;
wire n_10137;
wire n_10138;
wire n_10139;
wire n_10140;
wire n_10141;
wire n_10142;
wire n_10143;
wire n_10144;
wire n_10145;
wire n_10146;
wire n_10147;
wire n_10148;
wire n_10149;
wire n_10150;
wire n_10151;
wire n_10152;
wire n_10153;
wire n_10154;
wire n_10155;
wire n_10156;
wire n_10157;
wire n_10158;
wire n_10159;
wire n_10160;
wire n_10161;
wire n_10162;
wire n_10163;
wire n_10164;
wire n_10165;
wire n_10166;
wire n_10167;
wire n_10168;
wire n_10169;
wire n_10170;
wire n_10171;
wire n_10172;
wire n_10173;
wire n_10174;
wire n_10175;
wire n_10176;
wire n_10177;
wire n_10178;
wire n_10179;
wire n_10180;
wire n_10181;
wire n_10182;
wire n_10183;
wire n_10184;
wire n_10185;
wire n_10186;
wire n_10187;
wire n_10188;
wire n_10189;
wire n_10190;
wire n_10191;
wire n_10192;
wire n_10193;
wire n_10194;
wire n_10195;
wire n_10196;
wire n_10197;
wire n_10198;
wire n_10199;
wire n_10200;
wire n_10201;
wire n_10202;
wire n_10203;
wire n_10204;
wire n_10205;
wire n_10206;
wire n_10207;
wire n_10208;
wire n_10209;
wire n_10210;
wire n_10211;
wire n_10212;
wire n_10213;
wire n_10214;
wire n_10215;
wire n_10216;
wire n_10217;
wire n_10218;
wire n_10219;
wire n_10220;
wire n_10221;
wire n_10222;
wire n_10223;
wire n_10224;
wire n_10225;
wire n_10226;
wire n_10227;
wire n_10228;
wire n_10229;
wire n_10230;
wire n_10231;
wire n_10232;
wire n_10233;
wire n_10234;
wire n_10235;
wire n_10236;
wire n_10237;
wire n_10238;
wire n_10239;
wire n_10240;
wire n_10241;
wire n_10242;
wire n_10243;
wire n_10244;
wire n_10245;
wire n_10246;
wire n_10247;
wire n_10248;
wire n_10249;
wire n_10250;
wire n_10251;
wire n_10252;
wire n_10253;
wire n_10254;
wire n_10255;
wire n_10256;
wire n_10257;
wire n_10258;
wire n_10259;
wire n_10260;
wire n_10261;
wire n_10262;
wire n_10263;
wire n_10264;
wire n_10265;
wire n_10266;
wire n_10267;
wire n_10268;
wire n_10269;
wire n_10270;
wire n_10271;
wire n_10272;
wire n_10273;
wire n_10274;
wire n_10275;
wire n_10276;
wire n_10277;
wire n_10278;
wire n_10279;
wire n_10280;
wire n_10281;
wire n_10282;
wire n_10283;
wire n_10284;
wire n_10285;
wire n_10286;
wire n_10287;
wire n_10288;
wire n_10289;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10293;
wire n_10294;
wire n_10295;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10299;
wire n_10300;
wire n_10301;
wire n_10302;
wire n_10303;
wire n_10304;
wire n_10305;
wire n_10306;
wire n_10307;
wire n_10308;
wire n_10309;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10313;
wire n_10314;
wire n_10315;
wire n_10316;
wire n_10317;
wire n_10318;
wire n_10319;
wire n_10320;
wire n_10321;
wire n_10322;
wire n_10323;
wire n_10324;
wire n_10325;
wire n_10326;
wire n_10327;
wire n_10328;
wire n_10329;
wire n_10330;
wire n_10331;
wire n_10332;
wire n_10333;
wire n_10334;
wire n_10335;
wire n_10336;
wire n_10337;
wire n_10338;
wire n_10339;
wire n_10340;
wire n_10341;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10345;
wire n_10346;
wire n_10347;
wire n_10348;
wire n_10349;
wire n_10350;
wire n_10351;
wire n_10352;
wire n_10353;
wire n_10354;
wire n_10355;
wire n_10356;
wire n_10357;
wire n_10358;
wire n_10359;
wire n_10360;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10364;
wire n_10365;
wire n_10366;
wire n_10367;
wire n_10368;
wire n_10369;
wire n_10370;
wire n_10371;
wire n_10372;
wire n_10373;
wire n_10374;
wire n_10375;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_10379;
wire n_10380;
wire n_10381;
wire n_10382;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10387;
wire n_10388;
wire n_10389;
wire n_10390;
wire n_10391;
wire n_10392;
wire n_10393;
wire n_10394;
wire n_10395;
wire n_10396;
wire n_10397;
wire n_10398;
wire n_10399;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10403;
wire n_10404;
wire n_10405;
wire n_10406;
wire n_10407;
wire n_10408;
wire n_10409;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10415;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_10420;
wire n_10421;
wire n_10422;
wire n_10423;
wire n_10424;
wire n_10425;
wire n_10426;
wire n_10427;
wire n_10428;
wire n_10429;
wire n_10430;
wire n_10431;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10435;
wire n_10436;
wire n_10437;
wire n_10438;
wire n_10439;
wire n_10440;
wire n_10441;
wire n_10442;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10448;
wire n_10449;
wire n_10450;
wire n_10451;
wire n_10452;
wire n_10453;
wire n_10454;
wire n_10455;
wire n_10456;
wire n_10457;
wire n_10458;
wire n_10459;
wire n_10460;
wire n_10461;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10466;
wire n_10467;
wire n_10468;
wire n_10469;
wire n_10470;
wire n_10471;
wire n_10472;
wire n_10473;
wire n_10474;
wire n_10475;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_10480;
wire n_10481;
wire n_10482;
wire n_10483;
wire n_10484;
wire n_10485;
wire n_10486;
wire n_10487;
wire n_10488;
wire n_10489;
wire n_10490;
wire n_10491;
wire n_10492;
wire n_10493;
wire n_10494;
wire n_10495;
wire n_10496;
wire n_10497;
wire n_10498;
wire n_10499;
wire n_10500;
wire n_10501;
wire n_10502;
wire n_10503;
wire n_10504;
wire n_10505;
wire n_10506;
wire n_10507;
wire n_10508;
wire n_10509;
wire n_10510;
wire n_10511;
wire n_10512;
wire n_10513;
wire n_10514;
wire n_10515;
wire n_10516;
wire n_10517;
wire n_10518;
wire n_10519;
wire n_10520;
wire n_10521;
wire n_10522;
wire n_10523;
wire n_10524;
wire n_10525;
wire n_10526;
wire n_10527;
wire n_10528;
wire n_10529;
wire n_10530;
wire n_10531;
wire n_10532;
wire n_10533;
wire n_10534;
wire n_10535;
wire n_10536;
wire n_10537;
wire n_10538;
wire n_10539;
wire n_10540;
wire n_10541;
wire n_10542;
wire n_10543;
wire n_10544;
wire n_10545;
wire n_10546;
wire n_10547;
wire n_10548;
wire n_10549;
wire n_10550;
wire n_10551;
wire n_10552;
wire n_10553;
wire n_10554;
wire n_10555;
wire n_10556;
wire n_10557;
wire n_10558;
wire n_10559;
wire n_10560;
wire n_10561;
wire n_10562;
wire n_10563;
wire n_10564;
wire n_10565;
wire n_10566;
wire n_10567;
wire n_10568;
wire n_10569;
wire n_10570;
wire n_10571;
wire n_10572;
wire n_10573;
wire n_10574;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10578;
wire n_10579;
wire n_10580;
wire n_10581;
wire n_10582;
wire n_10583;
wire n_10584;
wire n_10585;
wire n_10586;
wire n_10587;
wire n_10588;
wire n_10589;
wire n_10590;
wire n_10591;
wire n_10592;
wire n_10593;
wire n_10594;
wire n_10595;
wire n_10596;
wire n_10597;
wire n_10598;
wire n_10599;
wire n_10600;
wire n_10601;
wire n_10602;
wire n_10603;
wire n_10604;
wire n_10605;
wire n_10606;
wire n_10607;
wire n_10608;
wire n_10609;
wire n_10610;
wire n_10611;
wire n_10612;
wire n_10613;
wire n_10614;
wire n_10615;
wire n_10616;
wire n_10617;
wire n_10618;
wire n_10619;
wire n_10620;
wire n_10621;
wire n_10622;
wire n_10623;
wire n_10624;
wire n_10625;
wire n_10626;
wire n_10627;
wire n_10628;
wire n_10629;
wire n_10630;
wire n_10631;
wire n_10632;
wire n_10633;
wire n_10634;
wire n_10635;
wire n_10636;
wire n_10637;
wire n_10638;
wire n_10639;
wire n_10640;
wire n_10641;
wire n_10642;
wire n_10643;
wire n_10644;
wire n_10645;
wire n_10646;
wire n_10647;
wire n_10648;
wire n_10649;
wire n_10650;
wire n_10651;
wire n_10652;
wire n_10653;
wire n_10654;
wire n_10655;
wire n_10656;
wire n_10657;
wire n_10658;
wire n_10659;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10663;
wire n_10664;
wire n_10665;
wire n_10666;
wire n_10667;
wire n_10668;
wire n_10669;
wire n_10670;
wire n_10671;
wire n_10672;
wire n_10673;
wire n_10674;
wire n_10675;
wire n_10676;
wire n_10677;
wire n_10678;
wire n_10679;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10683;
wire n_10684;
wire n_10685;
wire n_10686;
wire n_10687;
wire n_10688;
wire n_10689;
wire n_10690;
wire n_10691;
wire n_10692;
wire n_10693;
wire n_10694;
wire n_10695;
wire n_10696;
wire n_10697;
wire n_10698;
wire n_10699;
wire n_10700;
wire n_10701;
wire n_10702;
wire n_10703;
wire n_10704;
wire n_10705;
wire n_10706;
wire n_10707;
wire n_10708;
wire n_10709;
wire n_10710;
wire n_10711;
wire n_10712;
wire n_10713;
wire n_10714;
wire n_10715;
wire n_10716;
wire n_10717;
wire n_10718;
wire n_10719;
wire n_10720;
wire n_10721;
wire n_10722;
wire n_10723;
wire n_10724;
wire n_10725;
wire n_10726;
wire n_10727;
wire n_10728;
wire n_10729;
wire n_10730;
wire n_10731;
wire n_10732;
wire n_10733;
wire n_10734;
wire n_10735;
wire n_10736;
wire n_10737;
wire n_10738;
wire n_10739;
wire n_10740;
wire n_10741;
wire n_10742;
wire n_10743;
wire n_10744;
wire n_10745;
wire n_10746;
wire n_10747;
wire n_10748;
wire n_10749;
wire n_10750;
wire n_10751;
wire n_10752;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10756;
wire n_10757;
wire n_10758;
wire n_10759;
wire n_10760;
wire n_10761;
wire n_10762;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10766;
wire n_10767;
wire n_10768;
wire n_10769;
wire n_10770;
wire n_10771;
wire n_10772;
wire n_10773;
wire n_10774;
wire n_10775;
wire n_10776;
wire n_10777;
wire n_10778;
wire n_10779;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10783;
wire n_10784;
wire n_10785;
wire n_10786;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_10790;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10794;
wire n_10795;
wire n_10796;
wire n_10797;
wire n_10798;
wire n_10799;
wire n_10800;
wire n_10801;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10805;
wire n_10806;
wire n_10807;
wire n_10808;
wire n_10809;
wire n_10810;
wire n_10811;
wire n_10812;
wire n_10813;
wire n_10814;
wire n_10815;
wire n_10816;
wire n_10817;
wire n_10818;
wire n_10819;
wire n_10820;
wire n_10821;
wire n_10822;
wire n_10823;
wire n_10824;
wire n_10825;
wire n_10826;
wire n_10827;
wire n_10828;
wire n_10829;
wire n_10830;
wire n_10831;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10837;
wire n_10838;
wire n_10839;
wire n_10840;
wire n_10841;
wire n_10842;
wire n_10843;
wire n_10844;
wire n_10845;
wire n_10846;
wire n_10847;
wire n_10848;
wire n_10849;
wire n_10850;
wire n_10851;
wire n_10852;
wire n_10853;
wire n_10854;
wire n_10855;
wire n_10856;
wire n_10857;
wire n_10858;
wire n_10859;
wire n_10860;
wire n_10861;
wire n_10862;
wire n_10863;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10868;
wire n_10869;
wire n_10870;
wire n_10871;
wire n_10872;
wire n_10873;
wire n_10874;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_10878;
wire n_10879;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10883;
wire n_10884;
wire n_10885;
wire n_10886;
wire n_10887;
wire n_10888;
wire n_10889;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10893;
wire n_10894;
wire n_10895;
wire n_10896;
wire n_10897;
wire n_10898;
wire n_10899;
wire n_10900;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_10910;
wire n_10911;
wire n_10912;
wire n_10913;
wire n_10914;
wire n_10915;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_10920;
wire n_10921;
wire n_10922;
wire n_10923;
wire n_10924;
wire n_10925;
wire n_10926;
wire n_10927;
wire n_10928;
wire n_10929;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10933;
wire n_10934;
wire n_10935;
wire n_10936;
wire n_10937;
wire n_10938;
wire n_10939;
wire n_10940;
wire n_10941;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10945;
wire n_10946;
wire n_10947;
wire n_10948;
wire n_10949;
wire n_10950;
wire n_10951;
wire n_10952;
wire n_10953;
wire n_10954;
wire n_10955;
wire n_10956;
wire n_10957;
wire n_10958;
wire n_10959;
wire n_10960;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10964;
wire n_10965;
wire n_10966;
wire n_10967;
wire n_10968;
wire n_10969;
wire n_10970;
wire n_10971;
wire n_10972;
wire n_10973;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_10979;
wire n_10980;
wire n_10981;
wire n_10982;
wire n_10983;
wire n_10984;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_10988;
wire n_10989;
wire n_10990;
wire n_10991;
wire n_10992;
wire n_10993;
wire n_10994;
wire n_10995;
wire n_10996;
wire n_10997;
wire n_10998;
wire n_10999;
wire n_11000;
wire n_11001;
wire n_11002;
wire n_11003;
wire n_11004;
wire n_11005;
wire n_11006;
wire n_11007;
wire n_11008;
wire n_11009;
wire n_11010;
wire n_11011;
wire n_11012;
wire n_11013;
wire n_11014;
wire n_11015;
wire n_11016;
wire n_11017;
wire n_11018;
wire n_11019;
wire n_11020;
wire n_11021;
wire n_11022;
wire n_11023;
wire n_11024;
wire n_11025;
wire n_11026;
wire n_11027;
wire n_11028;
wire n_11029;
wire n_11030;
wire n_11031;
wire n_11032;
wire n_11033;
wire n_11034;
wire n_11035;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11045;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_11050;
wire n_11051;
wire n_11052;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11068;
wire n_11069;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11074;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_11080;
wire n_11081;
wire n_11082;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11098;
wire n_11099;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11103;
wire n_11104;
wire n_11105;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_11110;
wire n_11111;
wire n_11112;
wire n_11113;
wire n_11114;
wire n_11115;
wire n_11116;
wire n_11117;
wire n_11118;
wire n_11119;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11127;
wire n_11128;
wire n_11129;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11133;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_11140;
wire n_11141;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_11150;
wire n_11151;
wire n_11152;
wire n_11153;
wire n_11154;
wire n_11155;
wire n_11156;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_11160;
wire n_11161;
wire n_11162;
wire n_11163;
wire n_11164;
wire n_11165;
wire n_11166;
wire n_11167;
wire n_11168;
wire n_11169;
wire n_11170;
wire n_11171;
wire n_11172;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11176;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11183;
wire n_11184;
wire n_11185;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_11189;
wire n_11190;
wire n_11191;
wire n_11192;
wire n_11193;
wire n_11194;
wire n_11195;
wire n_11196;
wire n_11197;
wire n_11198;
wire n_11199;
wire n_11200;
wire n_11201;
wire n_11202;
wire n_11203;
wire n_11204;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_11210;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_11220;
wire n_11221;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11225;
wire n_11226;
wire n_11227;
wire n_11228;
wire n_11229;
wire n_11230;
wire n_11231;
wire n_11232;
wire n_11233;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11237;
wire n_11238;
wire n_11239;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11248;
wire n_11249;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11253;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11257;
wire n_11258;
wire n_11259;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11263;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11267;
wire n_11268;
wire n_11269;
wire n_11270;
wire n_11271;
wire n_11272;
wire n_11273;
wire n_11274;
wire n_11275;
wire n_11276;
wire n_11277;
wire n_11278;
wire n_11279;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11288;
wire n_11289;
wire n_11290;
wire n_11291;
wire n_11292;
wire n_11293;
wire n_11294;
wire n_11295;
wire n_11296;
wire n_11297;
wire n_11298;
wire n_11299;
wire n_11300;
wire n_11301;
wire n_11302;
wire n_11303;
wire n_11304;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11308;
wire n_11309;
wire n_11310;
wire n_11311;
wire n_11312;
wire n_11313;
wire n_11314;
wire n_11315;
wire n_11316;
wire n_11317;
wire n_11318;
wire n_11319;
wire n_11320;
wire n_11321;
wire n_11322;
wire n_11323;
wire n_11324;
wire n_11325;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_11329;
wire n_11330;
wire n_11331;
wire n_11332;
wire n_11333;
wire n_11334;
wire n_11335;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_11339;
wire n_11340;
wire n_11341;
wire n_11342;
wire n_11343;
wire n_11344;
wire n_11345;
wire n_11346;
wire n_11347;
wire n_11348;
wire n_11349;
wire n_11350;
wire n_11351;
wire n_11352;
wire n_11353;
wire n_11354;
wire n_11355;
wire n_11356;
wire n_11357;
wire n_11358;
wire n_11359;
wire n_11360;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11364;
wire n_11365;
wire n_11366;
wire n_11367;
wire n_11368;
wire n_11369;
wire n_11370;
wire n_11371;
wire n_11372;
wire n_11373;
wire n_11374;
wire n_11375;
wire n_11376;
wire n_11377;
wire n_11378;
wire n_11379;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11387;
wire n_11388;
wire n_11389;
wire n_11390;
wire n_11391;
wire n_11392;
wire n_11393;
wire n_11394;
wire n_11395;
wire n_11396;
wire n_11397;
wire n_11398;
wire n_11399;
wire n_11400;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11404;
wire n_11405;
wire n_11406;
wire n_11407;
wire n_11408;
wire n_11409;
wire n_11410;
wire n_11411;
wire n_11412;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11416;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_11420;
wire n_11421;
wire n_11422;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11426;
wire n_11427;
wire n_11428;
wire n_11429;
wire n_11430;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11439;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11444;
wire n_11445;
wire n_11446;
wire n_11447;
wire n_11448;
wire n_11449;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11453;
wire n_11454;
wire n_11455;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11459;
wire n_11460;
wire n_11461;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11465;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11469;
wire n_11470;
wire n_11471;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11475;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_11480;
wire n_11481;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11486;
wire n_11487;
wire n_11488;
wire n_11489;
wire n_11490;
wire n_11491;
wire n_11492;
wire n_11493;
wire n_11494;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11498;
wire n_11499;
wire n_11500;
wire n_11501;
wire n_11502;
wire n_11503;
wire n_11504;
wire n_11505;
wire n_11506;
wire n_11507;
wire n_11508;
wire n_11509;
wire n_11510;
wire n_11511;
wire n_11512;
wire n_11513;
wire n_11514;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11518;
wire n_11519;
wire n_11520;
wire n_11521;
wire n_11522;
wire n_11523;
wire n_11524;
wire n_11525;
wire n_11526;
wire n_11527;
wire n_11528;
wire n_11529;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11537;
wire n_11538;
wire n_11539;
wire n_11540;
wire n_11541;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_11550;
wire n_11551;
wire n_11552;
wire n_11553;
wire n_11554;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11558;
wire n_11559;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11563;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11567;
wire n_11568;
wire n_11569;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11574;
wire n_11575;
wire n_11576;
wire n_11577;
wire n_11578;
wire n_11579;
wire n_11580;
wire n_11581;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_11590;
wire n_11591;
wire n_11592;
wire n_11593;
wire n_11594;
wire n_11595;
wire n_11596;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11608;
wire n_11609;
wire n_11610;
wire n_11611;
wire n_11612;
wire n_11613;
wire n_11614;
wire n_11615;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_11619;
wire n_11620;
wire n_11621;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11627;
wire n_11628;
wire n_11629;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11636;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11643;
wire n_11644;
wire n_11645;
wire n_11646;
wire n_11647;
wire n_11648;
wire n_11649;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11654;
wire n_11655;
wire n_11656;
wire n_11657;
wire n_11658;
wire n_11659;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11664;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11673;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11678;
wire n_11679;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11704;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11709;
wire n_11710;
wire n_11711;
wire n_11712;
wire n_11713;
wire n_11714;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_11720;
wire n_11721;
wire n_11722;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_11729;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11737;
wire n_11738;
wire n_11739;
wire n_11740;
wire n_11741;
wire n_11742;
wire n_11743;
wire n_11744;
wire n_11745;
wire n_11746;
wire n_11747;
wire n_11748;
wire n_11749;
wire n_11750;
wire n_11751;
wire n_11752;
wire n_11753;
wire n_11754;
wire n_11755;
wire n_11756;
wire n_11757;
wire n_11758;
wire n_11759;
wire n_11760;
wire n_11761;
wire n_11762;
wire n_11763;
wire n_11764;
wire n_11765;
wire n_11766;
wire n_11767;
wire n_11768;
wire n_11769;
wire n_11770;
wire n_11771;
wire n_11772;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_11779;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11785;
wire n_11786;
wire n_11787;
wire n_11788;
wire n_11789;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11794;
wire n_11795;
wire n_11796;
wire n_11797;
wire n_11798;
wire n_11799;
wire n_11800;
wire n_11801;
wire n_11802;
wire n_11803;
wire n_11804;
wire n_11805;
wire n_11806;
wire n_11807;
wire n_11808;
wire n_11809;
wire n_11810;
wire n_11811;
wire n_11812;
wire n_11813;
wire n_11814;
wire n_11815;
wire n_11816;
wire n_11817;
wire n_11818;
wire n_11819;
wire n_11820;
wire n_11821;
wire n_11822;
wire n_11823;
wire n_11824;
wire n_11825;
wire n_11826;
wire n_11827;
wire n_11828;
wire n_11829;
wire n_11830;
wire n_11831;
wire n_11832;
wire n_11833;
wire n_11834;
wire n_11835;
wire n_11836;
wire n_11837;
wire n_11838;
wire n_11839;
wire n_11840;
wire n_11841;
wire n_11842;
wire n_11843;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_11879;
wire n_11880;
wire n_11881;
wire n_11882;
wire n_11883;
wire n_11884;
wire n_11885;
wire n_11886;
wire n_11887;
wire n_11888;
wire n_11889;
wire n_11890;
wire n_11891;
wire n_11892;
wire n_11893;
wire n_11894;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_11899;
wire n_11900;
wire n_11901;
wire n_11902;
wire n_11903;
wire n_11904;
wire n_11905;
wire n_11906;
wire n_11907;
wire n_11908;
wire n_11909;
wire n_11910;
wire n_11911;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire n_11916;
wire n_11917;
wire n_11918;
wire n_11919;
wire n_11920;
wire n_11921;
wire n_11922;
wire n_11923;
wire n_11924;
wire n_11925;
wire n_11926;
wire n_11927;
wire n_11928;
wire n_11929;
wire n_11930;
wire n_11931;
wire n_11932;
wire n_11933;
wire n_11934;
wire n_11935;
wire n_11936;
wire n_11937;
wire n_11938;
wire n_11939;
wire n_11940;
wire n_11941;
wire n_11942;
wire n_11943;
wire n_11944;
wire n_11945;
wire n_11946;
wire n_11947;
wire n_11948;
wire n_11949;
wire n_11950;
wire n_11951;
wire n_11952;
wire n_11953;
wire n_11954;
wire n_11955;
wire n_11956;
wire n_11957;
wire n_11958;
wire n_11959;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11963;
wire n_11964;
wire n_11965;
wire n_11966;
wire n_11967;
wire n_11968;
wire n_11969;
wire n_11970;
wire n_11971;
wire n_11972;
wire n_11973;
wire n_11974;
wire n_11975;
wire n_11976;
wire n_11977;
wire n_11978;
wire n_11979;
wire n_11980;
wire n_11981;
wire n_11982;
wire n_11983;
wire n_11984;
wire n_11985;
wire n_11986;
wire n_11987;
wire n_11988;
wire n_11989;
wire n_11990;
wire n_11991;
wire n_11992;
wire n_11993;
wire n_11994;
wire n_11995;
wire n_11996;
wire n_11997;
wire n_11998;
wire n_11999;
wire n_12000;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire n_12005;
wire n_12006;
wire n_12007;
wire n_12008;
wire n_12009;
wire n_12010;
wire n_12011;
wire n_12012;
wire n_12013;
wire n_12014;
wire n_12015;
wire n_12016;
wire n_12017;
wire n_12018;
wire n_12019;
wire n_12020;
wire n_12021;
wire n_12022;
wire n_12023;
wire n_12024;
wire n_12025;
wire n_12026;
wire n_12027;
wire n_12028;
wire n_12029;
wire n_12030;
wire n_12031;
wire n_12032;
wire n_12033;
wire n_12034;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_12039;
wire n_12040;
wire n_12041;
wire n_12042;
wire n_12043;
wire n_12044;
wire n_12045;
wire n_12046;
wire n_12047;
wire n_12048;
wire n_12049;
wire n_12050;
wire n_12051;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire n_12057;
wire n_12058;
wire n_12059;
wire n_12060;
wire n_12061;
wire n_12062;
wire n_12063;
wire n_12064;
wire n_12065;
wire n_12066;
wire n_12067;
wire n_12068;
wire n_12069;
wire n_12070;
wire n_12071;
wire n_12072;
wire n_12073;
wire n_12074;
wire n_12075;
wire n_12076;
wire n_12077;
wire n_12078;
wire n_12079;
wire n_12080;
wire n_12081;
wire n_12082;
wire n_12083;
wire n_12084;
wire n_12085;
wire n_12086;
wire n_12087;
wire n_12088;
wire n_12089;
wire n_12090;
wire n_12091;
wire n_12092;
wire n_12093;
wire n_12094;
wire n_12095;
wire n_12096;
wire n_12097;
wire n_12098;
wire n_12099;
wire n_12100;
wire n_12101;
wire n_12102;
wire n_12103;
wire n_12104;
wire n_12105;
wire n_12106;
wire n_12107;
wire n_12108;
wire n_12109;
wire n_12110;
wire n_12111;
wire n_12112;
wire n_12113;
wire n_12114;
wire n_12115;
wire n_12116;
wire n_12117;
wire n_12118;
wire n_12119;
wire n_12120;
wire n_12121;
wire n_12122;
wire n_12123;
wire n_12124;
wire n_12125;
wire n_12126;
wire n_12127;
wire n_12128;
wire n_12129;
wire n_12130;
wire n_12131;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12136;
wire n_12137;
wire n_12138;
wire n_12139;
wire n_12140;
wire n_12141;
wire n_12142;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_12149;
wire n_12150;
wire n_12151;
wire n_12152;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12157;
wire n_12158;
wire n_12159;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_12170;
wire n_12171;
wire n_12172;
wire n_12173;
wire n_12174;
wire n_12175;
wire n_12176;
wire n_12177;
wire n_12178;
wire n_12179;
wire n_12180;
wire n_12181;
wire n_12182;
wire n_12183;
wire n_12184;
wire n_12185;
wire n_12186;
wire n_12187;
wire n_12188;
wire n_12189;
wire n_12190;
wire n_12191;
wire n_12192;
wire n_12193;
wire n_12194;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire n_12199;
wire n_12200;
wire n_12201;
wire n_12202;
wire n_12203;
wire n_12204;
wire n_12205;
wire n_12206;
wire n_12207;
wire n_12208;
wire n_12209;
wire n_12210;
wire n_12211;
wire n_12212;
wire n_12213;
wire n_12214;
wire n_12215;
wire n_12216;
wire n_12217;
wire n_12218;
wire n_12219;
wire n_12220;
wire n_12221;
wire n_12222;
wire n_12223;
wire n_12224;
wire n_12225;
wire n_12226;
wire n_12227;
wire n_12228;
wire n_12229;
wire n_12230;
wire n_12231;
wire n_12232;
wire n_12233;
wire n_12234;
wire n_12235;
wire n_12236;
wire n_12237;
wire n_12238;
wire n_12239;
wire n_12240;
wire n_12241;
wire n_12242;
wire n_12243;
wire n_12244;
wire n_12245;
wire n_12246;
wire n_12247;
wire n_12248;
wire n_12249;
wire n_12250;
wire n_12251;
wire n_12252;
wire n_12253;
wire n_12254;
wire n_12255;
wire n_12256;
wire n_12257;
wire n_12258;
wire n_12259;
wire n_12260;
wire n_12261;
wire n_12262;
wire n_12263;
wire n_12264;
wire n_12265;
wire n_12266;
wire n_12267;
wire n_12268;
wire n_12269;
wire n_12270;
wire n_12271;
wire n_12272;
wire n_12273;
wire n_12274;
wire n_12275;
wire n_12276;
wire n_12277;
wire n_12278;
wire n_12279;
wire n_12280;
wire n_12281;
wire n_12282;
wire n_12283;
wire n_12284;
wire n_12285;
wire n_12286;
wire n_12287;
wire n_12288;
wire n_12289;
wire n_12290;
wire n_12291;
wire n_12292;
wire n_12293;
wire n_12294;
wire n_12295;
wire n_12296;
wire n_12297;
wire n_12298;
wire n_12299;
wire n_12300;
wire n_12301;
wire n_12302;
wire n_12303;
wire n_12304;
wire n_12305;
wire n_12306;
wire n_12307;
wire n_12308;
wire n_12309;
wire n_12310;
wire n_12311;
wire n_12312;
wire n_12313;
wire n_12314;
wire n_12315;
wire n_12316;
wire n_12317;
wire n_12318;
wire n_12319;
wire n_12320;
wire n_12321;
wire n_12322;
wire n_12323;
wire n_12324;
wire n_12325;
wire n_12326;
wire n_12327;
wire n_12328;
wire n_12329;
wire n_12330;
wire n_12331;
wire n_12332;
wire n_12333;
wire n_12334;
wire n_12335;
wire n_12336;
wire n_12337;
wire n_12338;
wire n_12339;
wire n_12340;
wire n_12341;
wire n_12342;
wire n_12343;
wire n_12344;
wire n_12345;
wire n_12346;
wire n_12347;
wire n_12348;
wire n_12349;
wire n_12350;
wire n_12351;
wire n_12352;
wire n_12353;
wire n_12354;
wire n_12355;
wire n_12356;
wire n_12357;
wire n_12358;
wire n_12359;
wire n_12360;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12364;
wire n_12365;
wire n_12366;
wire n_12367;
wire n_12368;
wire n_12369;
wire n_12370;
wire n_12371;
wire n_12372;
wire n_12373;
wire n_12374;
wire n_12375;
wire n_12376;
wire n_12377;
wire n_12378;
wire n_12379;
wire n_12380;
wire n_12381;
wire n_12382;
wire n_12383;
wire n_12384;
wire n_12385;
wire n_12386;
wire n_12387;
wire n_12388;
wire n_12389;
wire n_12390;
wire n_12391;
wire n_12392;
wire n_12393;
wire n_12394;
wire n_12395;
wire n_12396;
wire n_12397;
wire n_12398;
wire n_12399;
wire n_12400;
wire n_12401;
wire n_12402;
wire n_12403;
wire n_12404;
wire n_12405;
wire n_12406;
wire n_12407;
wire n_12408;
wire n_12409;
wire n_12410;
wire n_12411;
wire n_12412;
wire n_12413;
wire n_12414;
wire n_12415;
wire n_12416;
wire n_12417;
wire n_12418;
wire n_12419;
wire n_12420;
wire n_12421;
wire n_12422;
wire n_12423;
wire n_12424;
wire n_12425;
wire n_12426;
wire n_12427;
wire n_12428;
wire n_12429;
wire n_12430;
wire n_12431;
wire n_12432;
wire n_12433;
wire n_12434;
wire n_12435;
wire n_12436;
wire n_12437;
wire n_12438;
wire n_12439;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12443;
wire n_12444;
wire n_12445;
wire n_12446;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12456;
wire n_12457;
wire n_12458;
wire n_12459;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire n_12466;
wire n_12467;
wire n_12468;
wire n_12469;
wire n_12470;
wire n_12471;
wire n_12472;
wire n_12473;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12477;
wire n_12478;
wire n_12479;
wire n_12480;
wire n_12481;
wire n_12482;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12497;
wire n_12498;
wire n_12499;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12576;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_12580;
wire n_12581;
wire n_12582;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_12590;
wire n_12591;
wire n_12592;
wire n_12593;
wire n_12594;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_12600;
wire n_12601;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_12608;
wire n_12609;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12627;
wire n_12628;
wire n_12629;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12657;
wire n_12658;
wire n_12659;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12687;
wire n_12688;
wire n_12689;
wire n_12690;
wire n_12691;
wire n_12692;
wire n_12693;
wire n_12694;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12698;
wire n_12699;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12708;
wire n_12709;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_12718;
wire n_12719;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_12730;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_12739;
wire n_12740;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12755;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12777;
wire n_12778;
wire n_12779;
wire n_12780;
wire n_12781;
wire n_12782;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12793;
wire n_12794;
wire n_12795;
wire n_12796;
wire n_12797;
wire n_12798;
wire n_12799;
wire n_12800;
wire n_12801;
wire n_12802;
wire n_12803;
wire n_12804;
wire n_12805;
wire n_12806;
wire n_12807;
wire n_12808;
wire n_12809;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_12820;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12838;
wire n_12839;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12844;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12854;
wire n_12855;
wire n_12856;
wire n_12857;
wire n_12858;
wire n_12859;
wire n_12860;
wire n_12861;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_12909;
wire n_12910;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12925;
wire n_12926;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12944;
wire n_12945;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12953;
wire n_12954;
wire n_12955;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12965;
wire n_12966;
wire n_12967;
wire n_12968;
wire n_12969;
wire n_12970;
wire n_12971;
wire n_12972;
wire n_12973;
wire n_12974;
wire n_12975;
wire n_12976;
wire n_12977;
wire n_12978;
wire n_12979;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12987;
wire n_12988;
wire n_12989;
wire n_12990;
wire n_12991;
wire n_12992;
wire n_12993;
wire n_12994;
wire n_12995;
wire n_12996;
wire n_12997;
wire n_12998;
wire n_12999;
wire n_13000;
wire n_13001;
wire n_13002;
wire n_13003;
wire n_13004;
wire n_13005;
wire n_13006;
wire n_13007;
wire n_13008;
wire n_13009;
wire n_13010;
wire n_13011;
wire n_13012;
wire n_13013;
wire n_13014;
wire n_13015;
wire n_13016;
wire n_13017;
wire n_13018;
wire n_13019;
wire n_13020;
wire n_13021;
wire n_13022;
wire n_13023;
wire n_13024;
wire n_13025;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13029;
wire n_13030;
wire n_13031;
wire n_13032;
wire n_13033;
wire n_13034;
wire n_13035;
wire n_13036;
wire n_13037;
wire n_13038;
wire n_13039;
wire n_13040;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_13060;
wire n_13061;
wire n_13062;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13069;
wire n_13070;
wire n_13071;
wire n_13072;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_13090;
wire n_13091;
wire n_13092;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13096;
wire n_13097;
wire n_13098;
wire n_13099;
wire n_13100;
wire n_13101;
wire n_13102;
wire n_13103;
wire n_13104;
wire n_13105;
wire n_13106;
wire n_13107;
wire n_13108;
wire n_13109;
wire n_13110;
wire n_13111;
wire n_13112;
wire n_13113;
wire n_13114;
wire n_13115;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13119;
wire n_13120;
wire n_13121;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13126;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_13147;
wire n_13148;
wire n_13149;
wire n_13150;
wire n_13151;
wire n_13152;
wire n_13153;
wire n_13154;
wire n_13155;
wire n_13156;
wire n_13157;
wire n_13158;
wire n_13159;
wire n_13160;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_13169;
wire n_13170;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13174;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_13180;
wire n_13181;
wire n_13182;
wire n_13183;
wire n_13184;
wire n_13185;
wire n_13186;
wire n_13187;
wire n_13188;
wire n_13189;
wire n_13190;
wire n_13191;
wire n_13192;
wire n_13193;
wire n_13194;
wire n_13195;
wire n_13196;
wire n_13197;
wire n_13198;
wire n_13199;
wire n_13200;
wire n_13201;
wire n_13202;
wire n_13203;
wire n_13204;
wire n_13205;
wire n_13206;
wire n_13207;
wire n_13208;
wire n_13209;
wire n_13210;
wire n_13211;
wire n_13212;
wire n_13213;
wire n_13214;
wire n_13215;
wire n_13216;
wire n_13217;
wire n_13218;
wire n_13219;
wire n_13220;
wire n_13221;
wire n_13222;
wire n_13223;
wire n_13224;
wire n_13225;
wire n_13226;
wire n_13227;
wire n_13228;
wire n_13229;
wire n_13230;
wire n_13231;
wire n_13232;
wire n_13233;
wire n_13234;
wire n_13235;
wire n_13236;
wire n_13237;
wire n_13238;
wire n_13239;
wire n_13240;
wire n_13241;
wire n_13242;
wire n_13243;
wire n_13244;
wire n_13245;
wire n_13246;
wire n_13247;
wire n_13248;
wire n_13249;
wire n_13250;
wire n_13251;
wire n_13252;
wire n_13253;
wire n_13254;
wire n_13255;
wire n_13256;
wire n_13257;
wire n_13258;
wire n_13259;
wire n_13260;
wire n_13261;
wire n_13262;
wire n_13263;
wire n_13264;
wire n_13265;
wire n_13266;
wire n_13267;
wire n_13268;
wire n_13269;
wire n_13270;
wire n_13271;
wire n_13272;
wire n_13273;
wire n_13274;
wire n_13275;
wire n_13276;
wire n_13277;
wire n_13278;
wire n_13279;
wire n_13280;
wire n_13281;
wire n_13282;
wire n_13283;
wire n_13284;
wire n_13285;
wire n_13286;
wire n_13287;
wire n_13288;
wire n_13289;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13293;
wire n_13294;
wire n_13295;
wire n_13296;
wire n_13297;
wire n_13298;
wire n_13299;
wire n_13300;
wire n_13301;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13307;
wire n_13308;
wire n_13309;
wire n_13310;
wire n_13311;
wire n_13312;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13316;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_13320;
wire n_13321;
wire n_13322;
wire n_13323;
wire n_13324;
wire n_13325;
wire n_13326;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_13330;
wire n_13331;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire n_13336;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_13340;
wire n_13341;
wire n_13342;
wire n_13343;
wire n_13344;
wire n_13345;
wire n_13346;
wire n_13347;
wire n_13348;
wire n_13349;
wire n_13350;
wire n_13351;
wire n_13352;
wire n_13353;
wire n_13354;
wire n_13355;
wire n_13356;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13364;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_13380;
wire n_13381;
wire n_13382;
wire n_13383;
wire n_13384;
wire n_13385;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13396;
wire n_13397;
wire n_13398;
wire n_13399;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13413;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13433;
wire n_13434;
wire n_13435;
wire n_13436;
wire n_13437;
wire n_13438;
wire n_13439;
wire n_13440;
wire n_13441;
wire n_13442;
wire n_13443;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_13450;
wire n_13451;
wire n_13452;
wire n_13453;
wire n_13454;
wire n_13455;
wire n_13456;
wire n_13457;
wire n_13458;
wire n_13459;
wire n_13460;
wire n_13461;
wire n_13462;
wire n_13463;
wire n_13464;
wire n_13465;
wire n_13466;
wire n_13467;
wire n_13468;
wire n_13469;
wire n_13470;
wire n_13471;
wire n_13472;
wire n_13473;
wire n_13474;
wire n_13475;
wire n_13476;
wire n_13477;
wire n_13478;
wire n_13479;
wire n_13480;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire n_13489;
wire n_13490;
wire n_13491;
wire n_13492;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13498;
wire n_13499;
wire n_13500;
wire n_13501;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13507;
wire n_13508;
wire n_13509;
wire n_13510;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_13540;
wire n_13541;
wire n_13542;
wire n_13543;
wire n_13544;
wire n_13545;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_13549;
wire n_13550;
wire n_13551;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire n_13567;
wire n_13568;
wire n_13569;
wire n_13570;
wire n_13571;
wire n_13572;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_13580;
wire n_13581;
wire n_13582;
wire n_13583;
wire n_13584;
wire n_13585;
wire n_13586;
wire n_13587;
wire n_13588;
wire n_13589;
wire n_13590;
wire n_13591;
wire n_13592;
wire n_13593;
wire n_13594;
wire n_13595;
wire n_13596;
wire n_13597;
wire n_13598;
wire n_13599;
wire n_13600;
wire n_13601;
wire n_13602;
wire n_13603;
wire n_13604;
wire n_13605;
wire n_13606;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_13610;
wire n_13611;
wire n_13612;
wire n_13613;
wire n_13614;
wire n_13615;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13626;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_13630;
wire n_13631;
wire n_13632;
wire n_13633;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13637;
wire n_13638;
wire n_13639;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13644;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_13649;
wire n_13650;
wire n_13651;
wire n_13652;
wire n_13653;
wire n_13654;
wire n_13655;
wire n_13656;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_13660;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13665;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13669;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13675;
wire n_13676;
wire n_13677;
wire n_13678;
wire n_13679;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13683;
wire n_13684;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_13690;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13699;
wire n_13700;
wire n_13701;
wire n_13702;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13706;
wire n_13707;
wire n_13708;
wire n_13709;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13713;
wire n_13714;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13718;
wire n_13719;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13723;
wire n_13724;
wire n_13725;
wire n_13726;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_13730;
wire n_13731;
wire n_13732;
wire n_13733;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13737;
wire n_13738;
wire n_13739;
wire n_13740;
wire n_13741;
wire n_13742;
wire n_13743;
wire n_13744;
wire n_13745;
wire n_13746;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13751;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_13760;
wire n_13761;
wire n_13762;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_13769;
wire n_13770;
wire n_13771;
wire n_13772;
wire n_13773;
wire n_13774;
wire n_13775;
wire n_13776;
wire n_13777;
wire n_13778;
wire n_13779;
wire n_13780;
wire n_13781;
wire n_13782;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13786;
wire n_13787;
wire n_13788;
wire n_13789;
wire n_13790;
wire n_13791;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13795;
wire n_13796;
wire n_13797;
wire n_13798;
wire n_13799;
wire n_13800;
wire n_13801;
wire n_13802;
wire n_13803;
wire n_13804;
wire n_13805;
wire n_13806;
wire n_13807;
wire n_13808;
wire n_13809;
wire n_13810;
wire n_13811;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13818;
wire n_13819;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_13830;
wire n_13831;
wire n_13832;
wire n_13833;
wire n_13834;
wire n_13835;
wire n_13836;
wire n_13837;
wire n_13838;
wire n_13839;
wire n_13840;
wire n_13841;
wire n_13842;
wire n_13843;
wire n_13844;
wire n_13845;
wire n_13846;
wire n_13847;
wire n_13848;
wire n_13849;
wire n_13850;
wire n_13851;
wire n_13852;
wire n_13853;
wire n_13854;
wire n_13855;
wire n_13856;
wire n_13857;
wire n_13858;
wire n_13859;
wire n_13860;
wire n_13861;
wire n_13862;
wire n_13863;
wire n_13864;
wire n_13865;
wire n_13866;
wire n_13867;
wire n_13868;
wire n_13869;
wire n_13870;
wire n_13871;
wire n_13872;
wire n_13873;
wire n_13874;
wire n_13875;
wire n_13876;
wire n_13877;
wire n_13878;
wire n_13879;
wire n_13880;
wire n_13881;
wire n_13882;
wire n_13883;
wire n_13884;
wire n_13885;
wire n_13886;
wire n_13887;
wire n_13888;
wire n_13889;
wire n_13890;
wire n_13891;
wire n_13892;
wire n_13893;
wire n_13894;
wire n_13895;
wire n_13896;
wire n_13897;
wire n_13898;
wire n_13899;
wire n_13900;
wire n_13901;
wire n_13902;
wire n_13903;
wire n_13904;
wire n_13905;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_13909;
wire n_13910;
wire n_13911;
wire n_13912;
wire n_13913;
wire n_13914;
wire n_13915;
wire n_13916;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire n_13924;
wire n_13925;
wire n_13926;
wire n_13927;
wire n_13928;
wire n_13929;
wire n_13930;
wire n_13931;
wire n_13932;
wire n_13933;
wire n_13934;
wire n_13935;
wire n_13936;
wire n_13937;
wire n_13938;
wire n_13939;
wire n_13940;
wire n_13941;
wire n_13942;
wire n_13943;
wire n_13944;
wire n_13945;
wire n_13946;
wire n_13947;
wire n_13948;
wire n_13949;
wire n_13950;
wire n_13951;
wire n_13952;
wire n_13953;
wire n_13954;
wire n_13955;
wire n_13956;
wire n_13957;
wire n_13958;
wire n_13959;
wire n_13960;
wire n_13961;
wire n_13962;
wire n_13963;
wire n_13964;
wire n_13965;
wire n_13966;
wire n_13967;
wire n_13968;
wire n_13969;
wire n_13970;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire n_13975;
wire n_13976;
wire n_13977;
wire n_13978;
wire n_13979;
wire n_13980;
wire n_13981;
wire n_13982;
wire n_13983;
wire n_13984;
wire n_13985;
wire n_13986;
wire n_13987;
wire n_13988;
wire n_13989;
wire n_13990;
wire n_13991;
wire n_13992;
wire n_13993;
wire n_13994;
wire n_13995;
wire n_13996;
wire n_13997;
wire n_13998;
wire n_13999;
wire n_14000;
wire n_14001;
wire n_14002;
wire n_14003;
wire n_14004;
wire n_14005;
wire n_14006;
wire n_14007;
wire n_14008;
wire n_14009;
wire n_14010;
wire n_14011;
wire n_14012;
wire n_14013;
wire n_14014;
wire n_14015;
wire n_14016;
wire n_14017;
wire n_14018;
wire n_14019;
wire n_14020;
wire n_14021;
wire n_14022;
wire n_14023;
wire n_14024;
wire n_14025;
wire n_14026;
wire n_14027;
wire n_14028;
wire n_14029;
wire n_14030;
wire n_14031;
wire n_14032;
wire n_14033;
wire n_14034;
wire n_14035;
wire n_14036;
wire n_14037;
wire n_14038;
wire n_14039;
wire n_14040;
wire n_14041;
wire n_14042;
wire n_14043;
wire n_14044;
wire n_14045;
wire n_14046;
wire n_14047;
wire n_14048;
wire n_14049;
wire n_14050;
wire n_14051;
wire n_14052;
wire n_14053;
wire n_14054;
wire n_14055;
wire n_14056;
wire n_14057;
wire n_14058;
wire n_14059;
wire n_14060;
wire n_14061;
wire n_14062;
wire n_14063;
wire n_14064;
wire n_14065;
wire n_14066;
wire n_14067;
wire n_14068;
wire n_14069;
wire n_14070;
wire n_14071;
wire n_14072;
wire n_14073;
wire n_14074;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire n_14087;
wire n_14088;
wire n_14089;
wire n_14090;
wire n_14091;
wire n_14092;
wire n_14093;
wire n_14094;
wire n_14095;
wire n_14096;
wire n_14097;
wire n_14098;
wire n_14099;
wire n_14100;
wire n_14101;
wire n_14102;
wire n_14103;
wire n_14104;
wire n_14105;
wire n_14106;
wire n_14107;
wire n_14108;
wire n_14109;
wire n_14110;
wire n_14111;
wire n_14112;
wire n_14113;
wire n_14114;
wire n_14115;
wire n_14116;
wire n_14117;
wire n_14118;
wire n_14119;
wire n_14120;
wire n_14121;
wire n_14122;
wire n_14123;
wire n_14124;
wire n_14125;
wire n_14126;
wire n_14127;
wire n_14128;
wire n_14129;
wire n_14130;
wire n_14131;
wire n_14132;
wire n_14133;
wire n_14134;
wire n_14135;
wire n_14136;
wire n_14137;
wire n_14138;
wire n_14139;
wire n_14140;
wire n_14141;
wire n_14142;
wire n_14143;
wire n_14144;
wire n_14145;
wire n_14146;
wire n_14147;
wire n_14148;
wire n_14149;
wire n_14150;
wire n_14151;
wire n_14152;
wire n_14153;
wire n_14154;
wire n_14155;
wire n_14156;
wire n_14157;
wire n_14158;
wire n_14159;
wire n_14160;
wire n_14161;
wire n_14162;
wire n_14163;
wire n_14164;
wire n_14165;
wire n_14166;
wire n_14167;
wire n_14168;
wire n_14169;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14173;
wire n_14174;
wire n_14175;
wire n_14176;
wire n_14177;
wire n_14178;
wire n_14179;
wire n_14180;
wire n_14181;
wire n_14182;
wire n_14183;
wire n_14184;
wire n_14185;
wire n_14186;
wire n_14187;
wire n_14188;
wire n_14189;
wire n_14190;
wire n_14191;
wire n_14192;
wire n_14193;
wire n_14194;
wire n_14195;
wire n_14196;
wire n_14197;
wire n_14198;
wire n_14199;
wire n_14200;
wire n_14201;
wire n_14202;
wire n_14203;
wire n_14204;
wire n_14205;
wire n_14206;
wire n_14207;
wire n_14208;
wire n_14209;
wire n_14210;
wire n_14211;
wire n_14212;
wire n_14213;
wire n_14214;
wire n_14215;
wire n_14216;
wire n_14217;
wire n_14218;
wire n_14219;
wire n_14220;
wire n_14221;
wire n_14222;
wire n_14223;
wire n_14224;
wire n_14225;
wire n_14226;
wire n_14227;
wire n_14228;
wire n_14229;
wire n_14230;
wire n_14231;
wire n_14232;
wire n_14233;
wire n_14234;
wire n_14235;
wire n_14236;
wire n_14237;
wire n_14238;
wire n_14239;
wire n_14240;
wire n_14241;
wire n_14242;
wire n_14243;
wire n_14244;
wire n_14245;
wire n_14246;
wire n_14247;
wire n_14248;
wire n_14249;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_14259;
wire n_14260;
wire n_14261;
wire n_14262;
wire n_14263;
wire n_14264;
wire n_14265;
wire n_14266;
wire n_14267;
wire n_14268;
wire n_14269;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14276;
wire n_14277;
wire n_14278;
wire n_14279;
wire n_14280;
wire n_14281;
wire n_14282;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_14287;
wire n_14288;
wire n_14289;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14294;
wire n_14295;
wire n_14296;
wire n_14297;
wire n_14298;
wire n_14299;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14395;
wire n_14396;
wire n_14397;
wire n_14398;
wire n_14399;
wire n_14400;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14404;
wire n_14405;
wire n_14406;
wire n_14407;
wire n_14408;
wire n_14409;
wire n_14410;
wire n_14411;
wire n_14412;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14417;
wire n_14418;
wire n_14419;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14423;
wire n_14424;
wire n_14425;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_14450;
wire n_14451;
wire n_14452;
wire n_14453;
wire n_14454;
wire n_14455;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14463;
wire n_14464;
wire n_14465;
wire n_14466;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_14470;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14488;
wire n_14489;
wire n_14490;
wire n_14491;
wire n_14492;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14496;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_14500;
wire n_14501;
wire n_14502;
wire n_14503;
wire n_14504;
wire n_14505;
wire n_14506;
wire n_14507;
wire n_14508;
wire n_14509;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14516;
wire n_14517;
wire n_14518;
wire n_14519;
wire n_14520;
wire n_14521;
wire n_14522;
wire n_14523;
wire n_14524;
wire n_14525;
wire n_14526;
wire n_14527;
wire n_14528;
wire n_14529;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14533;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14537;
wire n_14538;
wire n_14539;
wire n_14540;
wire n_14541;
wire n_14542;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14546;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_14550;
wire n_14551;
wire n_14552;
wire n_14553;
wire n_14554;
wire n_14555;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_14560;
wire n_14561;
wire n_14562;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14568;
wire n_14569;
wire n_14570;
wire n_14571;
wire n_14572;
wire n_14573;
wire n_14574;
wire n_14575;
wire n_14576;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_14580;
wire n_14581;
wire n_14582;
wire n_14583;
wire n_14584;
wire n_14585;
wire n_14586;
wire n_14587;
wire n_14588;
wire n_14589;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_14600;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14606;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14647;
wire n_14648;
wire n_14649;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_14660;
wire n_14661;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_14670;
wire n_14671;
wire n_14672;
wire n_14673;
wire n_14674;
wire n_14675;
wire n_14676;
wire n_14677;
wire n_14678;
wire n_14679;
wire n_14680;
wire n_14681;
wire n_14682;
wire n_14683;
wire n_14684;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_14690;
wire n_14691;
wire n_14692;
wire n_14693;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14704;
wire n_14705;
wire n_14706;
wire n_14707;
wire n_14708;
wire n_14709;
wire n_14710;
wire n_14711;
wire n_14712;
wire n_14713;
wire n_14714;
wire n_14715;
wire n_14716;
wire n_14717;
wire n_14718;
wire n_14719;
wire n_14720;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14729;
wire n_14730;
wire n_14731;
wire n_14732;
wire n_14733;
wire n_14734;
wire n_14735;
wire n_14736;
wire n_14737;
wire n_14738;
wire n_14739;
wire n_14740;
wire n_14741;
wire n_14742;
wire n_14743;
wire n_14744;
wire n_14745;
wire n_14746;
wire n_14747;
wire n_14748;
wire n_14749;
wire n_14750;
wire n_14751;
wire n_14752;
wire n_14753;
wire n_14754;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14758;
wire n_14759;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_14770;
wire n_14771;
wire n_14772;
wire n_14773;
wire n_14774;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_14779;
wire n_14780;
wire n_14781;
wire n_14782;
wire n_14783;
wire n_14784;
wire n_14785;
wire n_14786;
wire n_14787;
wire n_14788;
wire n_14789;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14795;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_14800;
wire n_14801;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_14809;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_14820;
wire n_14821;
wire n_14822;
wire n_14823;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14827;
wire n_14828;
wire n_14829;
wire n_14830;
wire n_14831;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14835;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14843;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14857;
wire n_14858;
wire n_14859;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14868;
wire n_14869;
wire n_14870;
wire n_14871;
wire n_14872;
wire n_14873;
wire n_14874;
wire n_14875;
wire n_14876;
wire n_14877;
wire n_14878;
wire n_14879;
wire n_14880;
wire n_14881;
wire n_14882;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14886;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14935;
wire n_14936;
wire n_14937;
wire n_14938;
wire n_14939;
wire n_14940;
wire n_14941;
wire n_14942;
wire n_14943;
wire n_14944;
wire n_14945;
wire n_14946;
wire n_14947;
wire n_14948;
wire n_14949;
wire n_14950;
wire n_14951;
wire n_14952;
wire n_14953;
wire n_14954;
wire n_14955;
wire n_14956;
wire n_14957;
wire n_14958;
wire n_14959;
wire n_14960;
wire n_14961;
wire n_14962;
wire n_14963;
wire n_14964;
wire n_14965;
wire n_14966;
wire n_14967;
wire n_14968;
wire n_14969;
wire n_14970;
wire n_14971;
wire n_14972;
wire n_14973;
wire n_14974;
wire n_14975;
wire n_14976;
wire n_14977;
wire n_14978;
wire n_14979;
wire n_14980;
wire n_14981;
wire n_14982;
wire n_14983;
wire n_14984;
wire n_14985;
wire n_14986;
wire n_14987;
wire n_14988;
wire n_14989;
wire n_14990;
wire n_14991;
wire n_14992;
wire n_14993;
wire n_14994;
wire n_14995;
wire n_14996;
wire n_14997;
wire n_14998;
wire n_14999;
wire n_15000;
wire n_15001;
wire n_15002;
wire n_15003;
wire n_15004;
wire n_15005;
wire n_15006;
wire n_15007;
wire n_15008;
wire n_15009;
wire n_15010;
wire n_15011;
wire n_15012;
wire n_15013;
wire n_15014;
wire n_15015;
wire n_15016;
wire n_15017;
wire n_15018;
wire n_15019;
wire n_15020;
wire n_15021;
wire n_15022;
wire n_15023;
wire n_15024;
wire n_15025;
wire n_15026;
wire n_15027;
wire n_15028;
wire n_15029;
wire n_15030;
wire n_15031;
wire n_15032;
wire n_15033;
wire n_15034;
wire n_15035;
wire n_15036;
wire n_15037;
wire n_15038;
wire n_15039;
wire n_15040;
wire n_15041;
wire n_15042;
wire n_15043;
wire n_15044;
wire n_15045;
wire n_15046;
wire n_15047;
wire n_15048;
wire n_15049;
wire n_15050;
wire n_15051;
wire n_15052;
wire n_15053;
wire n_15054;
wire n_15055;
wire n_15056;
wire n_15057;
wire n_15058;
wire n_15059;
wire n_15060;
wire n_15061;
wire n_15062;
wire n_15063;
wire n_15064;
wire n_15065;
wire n_15066;
wire n_15067;
wire n_15068;
wire n_15069;
wire n_15070;
wire n_15071;
wire n_15072;
wire n_15073;
wire n_15074;
wire n_15075;
wire n_15076;
wire n_15077;
wire n_15078;
wire n_15079;
wire n_15080;
wire n_15081;
wire n_15082;
wire n_15083;
wire n_15084;
wire n_15085;
wire n_15086;
wire n_15087;
wire n_15088;
wire n_15089;
wire n_15090;
wire n_15091;
wire n_15092;
wire n_15093;
wire n_15094;
wire n_15095;
wire n_15096;
wire n_15097;
wire n_15098;
wire n_15099;
wire n_15100;
wire n_15101;
wire n_15102;
wire n_15103;
wire n_15104;
wire n_15105;
wire n_15106;
wire n_15107;
wire n_15108;
wire n_15109;
wire n_15110;
wire n_15111;
wire n_15112;
wire n_15113;
wire n_15114;
wire n_15115;
wire n_15116;
wire n_15117;
wire n_15118;
wire n_15119;
wire n_15120;
wire n_15121;
wire n_15122;
wire n_15123;
wire n_15124;
wire n_15125;
wire n_15126;
wire n_15127;
wire n_15128;
wire n_15129;
wire n_15130;
wire n_15131;
wire n_15132;
wire n_15133;
wire n_15134;
wire n_15135;
wire n_15136;
wire n_15137;
wire n_15138;
wire n_15139;
wire n_15140;
wire n_15141;
wire n_15142;
wire n_15143;
wire n_15144;
wire n_15145;
wire n_15146;
wire n_15147;
wire n_15148;
wire n_15149;
wire n_15150;
wire n_15151;
wire n_15152;
wire n_15153;
wire n_15154;
wire n_15155;
wire n_15156;
wire n_15157;
wire n_15158;
wire n_15159;
wire n_15160;
wire n_15161;
wire n_15162;
wire n_15163;
wire n_15164;
wire n_15165;
wire n_15166;
wire n_15167;
wire n_15168;
wire n_15169;
wire n_15170;
wire n_15171;
wire n_15172;
wire n_15173;
wire n_15174;
wire n_15175;
wire n_15176;
wire n_15177;
wire n_15178;
wire n_15179;
wire n_15180;
wire n_15181;
wire n_15182;
wire n_15183;
wire n_15184;
wire n_15185;
wire n_15186;
wire n_15187;
wire n_15188;
wire n_15189;
wire n_15190;
wire n_15191;
wire n_15192;
wire n_15193;
wire n_15194;
wire n_15195;
wire n_15196;
wire n_15197;
wire n_15198;
wire n_15199;
wire n_15200;
wire n_15201;
wire n_15202;
wire n_15203;
wire n_15204;
wire n_15205;
wire n_15206;
wire n_15207;
wire n_15208;
wire n_15209;
wire n_15210;
wire n_15211;
wire n_15212;
wire n_15213;
wire n_15214;
wire n_15215;
wire n_15216;
wire n_15217;
wire n_15218;
wire n_15219;
wire n_15220;
wire n_15221;
wire n_15222;
wire n_15223;
wire n_15224;
wire n_15225;
wire n_15226;
wire n_15227;
wire n_15228;
wire n_15229;
wire n_15230;
wire n_15231;
wire n_15232;
wire n_15233;
wire n_15234;
wire n_15235;
wire n_15236;
wire n_15237;
wire n_15238;
wire n_15239;
wire n_15240;
wire n_15241;
wire n_15242;
wire n_15243;
wire n_15244;
wire n_15245;
wire n_15246;
wire n_15247;
wire n_15248;
wire n_15249;
wire n_15250;
wire n_15251;
wire n_15252;
wire n_15253;
wire n_15254;
wire n_15255;
wire n_15256;
wire n_15257;
wire n_15258;
wire n_15259;
wire n_15260;
wire n_15261;
wire n_15262;
wire n_15263;
wire n_15264;
wire n_15265;
wire n_15266;
wire n_15267;
wire n_15268;
wire n_15269;
wire n_15270;
wire n_15271;
wire n_15272;
wire n_15273;
wire n_15274;
wire n_15275;
wire n_15276;
wire n_15277;
wire n_15278;
wire n_15279;
wire n_15280;
wire n_15281;
wire n_15282;
wire n_15283;
wire n_15284;
wire n_15285;
wire n_15286;
wire n_15287;
wire n_15288;
wire n_15289;
wire n_15290;
wire n_15291;
wire n_15292;
wire n_15293;
wire n_15294;
wire n_15295;
wire n_15296;
wire n_15297;
wire n_15298;
wire n_15299;
wire n_15300;
wire n_15301;
wire n_15302;
wire n_15303;
wire n_15304;
wire n_15305;
wire n_15306;
wire n_15307;
wire n_15308;
wire n_15309;
wire n_15310;
wire n_15311;
wire n_15312;
wire n_15313;
wire n_15314;
wire n_15315;
wire n_15316;
wire n_15317;
wire n_15318;
wire n_15319;
wire n_15320;
wire n_15321;
wire n_15322;
wire n_15323;
wire n_15324;
wire n_15325;
wire n_15326;
wire n_15327;
wire n_15328;
wire n_15329;
wire n_15330;
wire n_15331;
wire n_15332;
wire n_15333;
wire n_15334;
wire n_15335;
wire n_15336;
wire n_15337;
wire n_15338;
wire n_15339;
wire n_15340;
wire n_15341;
wire n_15342;
wire n_15343;
wire n_15344;
wire n_15345;
wire n_15346;
wire n_15347;
wire n_15348;
wire n_15349;
wire n_15350;
wire n_15351;
wire n_15352;
wire n_15353;
wire n_15354;
wire n_15355;
wire n_15356;
wire n_15357;
wire n_15358;
wire n_15359;
wire n_15360;
wire n_15361;
wire n_15362;
wire n_15363;
wire n_15364;
wire n_15365;
wire n_15366;
wire n_15367;
wire n_15368;
wire n_15369;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15374;
wire n_15375;
wire n_15376;
wire n_15377;
wire n_15378;
wire n_15379;
wire n_15380;
wire n_15381;
wire n_15382;
wire n_15383;
wire n_15384;
wire n_15385;
wire n_15386;
wire n_15387;
wire n_15388;
wire n_15389;
wire n_15390;
wire n_15391;
wire n_15392;
wire n_15393;
wire n_15394;
wire n_15395;
wire n_15396;
wire n_15397;
wire n_15398;
wire n_15399;
wire n_15400;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15404;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_15408;
wire n_15409;
wire n_15410;
wire n_15411;
wire n_15412;
wire n_15413;
wire n_15414;
wire n_15415;
wire n_15416;
wire n_15417;
wire n_15418;
wire n_15419;
wire n_15420;
wire n_15421;
wire n_15422;
wire n_15423;
wire n_15424;
wire n_15425;
wire n_15426;
wire n_15427;
wire n_15428;
wire n_15429;
wire n_15430;
wire n_15431;
wire n_15432;
wire n_15433;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15437;
wire n_15438;
wire n_15439;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15443;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_15447;
wire n_15448;
wire n_15449;
wire n_15450;
wire n_15451;
wire n_15452;
wire n_15453;
wire n_15454;
wire n_15455;
wire n_15456;
wire n_15457;
wire n_15458;
wire n_15459;
wire n_15460;
wire n_15461;
wire n_15462;
wire n_15463;
wire n_15464;
wire n_15465;
wire n_15466;
wire n_15467;
wire n_15468;
wire n_15469;
wire n_15470;
wire n_15471;
wire n_15472;
wire n_15473;
wire n_15474;
wire n_15475;
wire n_15476;
wire n_15477;
wire n_15478;
wire n_15479;
wire n_15480;
wire n_15481;
wire n_15482;
wire n_15483;
wire n_15484;
wire n_15485;
wire n_15486;
wire n_15487;
wire n_15488;
wire n_15489;
wire n_15490;
wire n_15491;
wire n_15492;
wire n_15493;
wire n_15494;
wire n_15495;
wire n_15496;
wire n_15497;
wire n_15498;
wire n_15499;
wire n_15500;
wire n_15501;
wire n_15502;
wire n_15503;
wire n_15504;
wire n_15505;
wire n_15506;
wire n_15507;
wire n_15508;
wire n_15509;
wire n_15510;
wire n_15511;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire n_15519;
wire n_15520;
wire n_15521;
wire n_15522;
wire n_15523;
wire n_15524;
wire n_15525;
wire n_15526;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_15530;
wire n_15531;
wire n_15532;
wire n_15533;
wire n_15534;
wire n_15535;
wire n_15536;
wire n_15537;
wire n_15538;
wire n_15539;
wire n_15540;
wire n_15541;
wire n_15542;
wire n_15543;
wire n_15544;
wire n_15545;
wire n_15546;
wire n_15547;
wire n_15548;
wire n_15549;
wire n_15550;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15554;
wire n_15555;
wire n_15556;
wire n_15557;
wire n_15558;
wire n_15559;
wire n_15560;
wire n_15561;
wire n_15562;
wire n_15563;
wire n_15564;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_15570;
wire n_15571;
wire n_15572;
wire n_15573;
wire n_15574;
wire n_15575;
wire n_15576;
wire n_15577;
wire n_15578;
wire n_15579;
wire n_15580;
wire n_15581;
wire n_15582;
wire n_15583;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15588;
wire n_15589;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15595;
wire n_15596;
wire n_15597;
wire n_15598;
wire n_15599;
wire n_15600;
wire n_15601;
wire n_15602;
wire n_15603;
wire n_15604;
wire n_15605;
wire n_15606;
wire n_15607;
wire n_15608;
wire n_15609;
wire n_15610;
wire n_15611;
wire n_15612;
wire n_15613;
wire n_15614;
wire n_15615;
wire n_15616;
wire n_15617;
wire n_15618;
wire n_15619;
wire n_15620;
wire n_15621;
wire n_15622;
wire n_15623;
wire n_15624;
wire n_15625;
wire n_15626;
wire n_15627;
wire n_15628;
wire n_15629;
wire n_15630;
wire n_15631;
wire n_15632;
wire n_15633;
wire n_15634;
wire n_15635;
wire n_15636;
wire n_15637;
wire n_15638;
wire n_15639;
wire n_15640;
wire n_15641;
wire n_15642;
wire n_15643;
wire n_15644;
wire n_15645;
wire n_15646;
wire n_15647;
wire n_15648;
wire n_15649;
wire n_15650;
wire n_15651;
wire n_15652;
wire n_15653;
wire n_15654;
wire n_15655;
wire n_15656;
wire n_15657;
wire n_15658;
wire n_15659;
wire n_15660;
wire n_15661;
wire n_15662;
wire n_15663;
wire n_15664;
wire n_15665;
wire n_15666;
wire n_15667;
wire n_15668;
wire n_15669;
wire n_15670;
wire n_15671;
wire n_15672;
wire n_15673;
wire n_15674;
wire n_15675;
wire n_15676;
wire n_15677;
wire n_15678;
wire n_15679;
wire n_15680;
wire n_15681;
wire n_15682;
wire n_15683;
wire n_15684;
wire n_15685;
wire n_15686;
wire n_15687;
wire n_15688;
wire n_15689;
wire n_15690;
wire n_15691;
wire n_15692;
wire n_15693;
wire n_15694;
wire n_15695;
wire n_15696;
wire n_15697;
wire n_15698;
wire n_15699;
wire n_15700;
wire n_15701;
wire n_15702;
wire n_15703;
wire n_15704;
wire n_15705;
wire n_15706;
wire n_15707;
wire n_15708;
wire n_15709;
wire n_15710;
wire n_15711;
wire n_15712;
wire n_15713;
wire n_15714;
wire n_15715;
wire n_15716;
wire n_15717;
wire n_15718;
wire n_15719;
wire n_15720;
wire n_15721;
wire n_15722;
wire n_15723;
wire n_15724;
wire n_15725;
wire n_15726;
wire n_15727;
wire n_15728;
wire n_15729;
wire n_15730;
wire n_15731;
wire n_15732;
wire n_15733;
wire n_15734;
wire n_15735;
wire n_15736;
wire n_15737;
wire n_15738;
wire n_15739;
wire n_15740;
wire n_15741;
wire n_15742;
wire n_15743;
wire n_15744;
wire n_15745;
wire n_15746;
wire n_15747;
wire n_15748;
wire n_15749;
wire n_15750;
wire n_15751;
wire n_15752;
wire n_15753;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire n_15760;
wire n_15761;
wire n_15762;
wire n_15763;
wire n_15764;
wire n_15765;
wire n_15766;
wire n_15767;
wire n_15768;
wire n_15769;
wire n_15770;
wire n_15771;
wire n_15772;
wire n_15773;
wire n_15774;
wire n_15775;
wire n_15776;
wire n_15777;
wire n_15778;
wire n_15779;
wire n_15780;
wire n_15781;
wire n_15782;
wire n_15783;
wire n_15784;
wire n_15785;
wire n_15786;
wire n_15787;
wire n_15788;
wire n_15789;
wire n_15790;
wire n_15791;
wire n_15792;
wire n_15793;
wire n_15794;
wire n_15795;
wire n_15796;
wire n_15797;
wire n_15798;
wire n_15799;
wire n_15800;
wire n_15801;
wire n_15802;
wire n_15803;
wire n_15804;
wire n_15805;
wire n_15806;
wire n_15807;
wire n_15808;
wire n_15809;
wire n_15810;
wire n_15811;
wire n_15812;
wire n_15813;
wire n_15814;
wire n_15815;
wire n_15816;
wire n_15817;
wire n_15818;
wire n_15819;
wire n_15820;
wire n_15821;
wire n_15822;
wire n_15823;
wire n_15824;
wire n_15825;
wire n_15826;
wire n_15827;
wire n_15828;
wire n_15829;
wire n_15830;
wire n_15831;
wire n_15832;
wire n_15833;
wire n_15834;
wire n_15835;
wire n_15836;
wire n_15837;
wire n_15838;
wire n_15839;
wire n_15840;
wire n_15841;
wire n_15842;
wire n_15843;
wire n_15844;
wire n_15845;
wire n_15846;
wire n_15847;
wire n_15848;
wire n_15849;
wire n_15850;
wire n_15851;
wire n_15852;
wire n_15853;
wire n_15854;
wire n_15855;
wire n_15856;
wire n_15857;
wire n_15858;
wire n_15859;
wire n_15860;
wire n_15861;
wire n_15862;
wire n_15863;
wire n_15864;
wire n_15865;
wire n_15866;
wire n_15867;
wire n_15868;
wire n_15869;
wire n_15870;
wire n_15871;
wire n_15872;
wire n_15873;
wire n_15874;
wire n_15875;
wire n_15876;
wire n_15877;
wire n_15878;
wire n_15879;
wire n_15880;
wire n_15881;
wire n_15882;
wire n_15883;
wire n_15884;
wire n_15885;
wire n_15886;
wire n_15887;
wire n_15888;
wire n_15889;
wire n_15890;
wire n_15891;
wire n_15892;
wire n_15893;
wire n_15894;
wire n_15895;
wire n_15896;
wire n_15897;
wire n_15898;
wire n_15899;
wire n_15900;
wire n_15901;
wire n_15902;
wire n_15903;
wire n_15904;
wire n_15905;
wire n_15906;
wire n_15907;
wire n_15908;
wire n_15909;
wire n_15910;
wire n_15911;
wire n_15912;
wire n_15913;
wire n_15914;
wire n_15915;
wire n_15916;
wire n_15917;
wire n_15918;
wire n_15919;
wire n_15920;
wire n_15921;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15925;
wire n_15926;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_15930;
wire n_15931;
wire n_15932;
wire n_15933;
wire n_15934;
wire n_15935;
wire n_15936;
wire n_15937;
wire n_15938;
wire n_15939;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_15943;
wire n_15944;
wire n_15945;
wire n_15946;
wire n_15947;
wire n_15948;
wire n_15949;
wire n_15950;
wire n_15951;
wire n_15952;
wire n_15953;
wire n_15954;
wire n_15955;
wire n_15956;
wire n_15957;
wire n_15958;
wire n_15959;
wire n_15960;
wire n_15961;
wire n_15962;
wire n_15963;
wire n_15964;
wire n_15965;
wire n_15966;
wire n_15967;
wire n_15968;
wire n_15969;
wire n_15970;
wire n_15971;
wire n_15972;
wire n_15973;
wire n_15974;
wire n_15975;
wire n_15976;
wire n_15977;
wire n_15978;
wire n_15979;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15983;
wire n_15984;
wire n_15985;
wire n_15986;
wire n_15987;
wire n_15988;
wire n_15989;
wire n_15990;
wire n_15991;
wire n_15992;
wire n_15993;
wire n_15994;
wire n_15995;
wire n_15996;
wire n_15997;
wire n_15998;
wire n_15999;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_16004;
wire n_16005;
wire n_16006;
wire n_16007;
wire n_16008;
wire n_16009;
wire n_16010;
wire n_16011;
wire n_16012;
wire n_16013;
wire n_16014;
wire n_16015;
wire n_16016;
wire n_16017;
wire n_16018;
wire n_16019;
wire n_16020;
wire n_16021;
wire n_16022;
wire n_16023;
wire n_16024;
wire n_16025;
wire n_16026;
wire n_16027;
wire n_16028;
wire n_16029;
wire n_16030;
wire n_16031;
wire n_16032;
wire n_16033;
wire n_16034;
wire n_16035;
wire n_16036;
wire n_16037;
wire n_16038;
wire n_16039;
wire n_16040;
wire n_16041;
wire n_16042;
wire n_16043;
wire n_16044;
wire n_16045;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_16050;
wire n_16051;
wire n_16052;
wire n_16053;
wire n_16054;
wire n_16055;
wire n_16056;
wire n_16057;
wire n_16058;
wire n_16059;
wire n_16060;
wire n_16061;
wire n_16062;
wire n_16063;
wire n_16064;
wire n_16065;
wire n_16066;
wire n_16067;
wire n_16068;
wire n_16069;
wire n_16070;
wire n_16071;
wire n_16072;
wire n_16073;
wire n_16074;
wire n_16075;
wire n_16076;
wire n_16077;
wire n_16078;
wire n_16079;
wire n_16080;
wire n_16081;
wire n_16082;
wire n_16083;
wire n_16084;
wire n_16085;
wire n_16086;
wire n_16087;
wire n_16088;
wire n_16089;
wire n_16090;
wire n_16091;
wire n_16092;
wire n_16093;
wire n_16094;
wire n_16095;
wire n_16096;
wire n_16097;
wire n_16098;
wire n_16099;
wire n_16100;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16104;
wire n_16105;
wire n_16106;
wire n_16107;
wire n_16108;
wire n_16109;
wire n_16110;
wire n_16111;
wire n_16112;
wire n_16113;
wire n_16114;
wire n_16115;
wire n_16116;
wire n_16117;
wire n_16118;
wire n_16119;
wire n_16120;
wire n_16121;
wire n_16122;
wire n_16123;
wire n_16124;
wire n_16125;
wire n_16126;
wire n_16127;
wire n_16128;
wire n_16129;
wire n_16130;
wire n_16131;
wire n_16132;
wire n_16133;
wire n_16134;
wire n_16135;
wire n_16136;
wire n_16137;
wire n_16138;
wire n_16139;
wire n_16140;
wire n_16141;
wire n_16142;
wire n_16143;
wire n_16144;
wire n_16145;
wire n_16146;
wire n_16147;
wire n_16148;
wire n_16149;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16155;
wire n_16156;
wire n_16157;
wire n_16158;
wire n_16159;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire n_16166;
wire n_16167;
wire n_16168;
wire n_16169;
wire n_16170;
wire n_16171;
wire n_16172;
wire n_16173;
wire n_16174;
wire n_16175;
wire n_16176;
wire n_16177;
wire n_16178;
wire n_16179;
wire n_16180;
wire n_16181;
wire n_16182;
wire n_16183;
wire n_16184;
wire n_16185;
wire n_16186;
wire n_16187;
wire n_16188;
wire n_16189;
wire n_16190;
wire n_16191;
wire n_16192;
wire n_16193;
wire n_16194;
wire n_16195;
wire n_16196;
wire n_16197;
wire n_16198;
wire n_16199;
wire n_16200;
wire n_16201;
wire n_16202;
wire n_16203;
wire n_16204;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16214;
wire n_16215;
wire n_16216;
wire n_16217;
wire n_16218;
wire n_16219;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_16230;
wire n_16231;
wire n_16232;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_16240;
wire n_16241;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16245;
wire n_16246;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16263;
wire n_16264;
wire n_16265;
wire n_16266;
wire n_16267;
wire n_16268;
wire n_16269;
wire n_16270;
wire n_16271;
wire n_16272;
wire n_16273;
wire n_16274;
wire n_16275;
wire n_16276;
wire n_16277;
wire n_16278;
wire n_16279;
wire n_16280;
wire n_16281;
wire n_16282;
wire n_16283;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_16290;
wire n_16291;
wire n_16292;
wire n_16293;
wire n_16294;
wire n_16295;
wire n_16296;
wire n_16297;
wire n_16298;
wire n_16299;
wire n_16300;
wire n_16301;
wire n_16302;
wire n_16303;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16308;
wire n_16309;
wire n_16310;
wire n_16311;
wire n_16312;
wire n_16313;
wire n_16314;
wire n_16315;
wire n_16316;
wire n_16317;
wire n_16318;
wire n_16319;
wire n_16320;
wire n_16321;
wire n_16322;
wire n_16323;
wire n_16324;
wire n_16325;
wire n_16326;
wire n_16327;
wire n_16328;
wire n_16329;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16333;
wire n_16334;
wire n_16335;
wire n_16336;
wire n_16337;
wire n_16338;
wire n_16339;
wire n_16340;
wire n_16341;
wire n_16342;
wire n_16343;
wire n_16344;
wire n_16345;
wire n_16346;
wire n_16347;
wire n_16348;
wire n_16349;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16353;
wire n_16354;
wire n_16355;
wire n_16356;
wire n_16357;
wire n_16358;
wire n_16359;
wire n_16360;
wire n_16361;
wire n_16362;
wire n_16363;
wire n_16364;
wire n_16365;
wire n_16366;
wire n_16367;
wire n_16368;
wire n_16369;
wire n_16370;
wire n_16371;
wire n_16372;
wire n_16373;
wire n_16374;
wire n_16375;
wire n_16376;
wire n_16377;
wire n_16378;
wire n_16379;
wire n_16380;
wire n_16381;
wire n_16382;
wire n_16383;
wire n_16384;
wire n_16385;
wire n_16386;
wire n_16387;
wire n_16388;
wire n_16389;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16393;
wire n_16394;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16405;
wire n_16406;
wire n_16407;
wire n_16408;
wire n_16409;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_16414;
wire n_16415;
wire n_16416;
wire n_16417;
wire n_16418;
wire n_16419;
wire n_16420;
wire n_16421;
wire n_16422;
wire n_16423;
wire n_16424;
wire n_16425;
wire n_16426;
wire n_16427;
wire n_16428;
wire n_16429;
wire n_16430;
wire n_16431;
wire n_16432;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_16440;
wire n_16441;
wire n_16442;
wire n_16443;
wire n_16444;
wire n_16445;
wire n_16446;
wire n_16447;
wire n_16448;
wire n_16449;
wire n_16450;
wire n_16451;
wire n_16452;
wire n_16453;
wire n_16454;
wire n_16455;
wire n_16456;
wire n_16457;
wire n_16458;
wire n_16459;
wire n_16460;
wire n_16461;
wire n_16462;
wire n_16463;
wire n_16464;
wire n_16465;
wire n_16466;
wire n_16467;
wire n_16468;
wire n_16469;
wire n_16470;
wire n_16471;
wire n_16472;
wire n_16473;
wire n_16474;
wire n_16475;
wire n_16476;
wire n_16477;
wire n_16478;
wire n_16479;
wire n_16480;
wire n_16481;
wire n_16482;
wire n_16483;
wire n_16484;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_16488;
wire n_16489;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16498;
wire n_16499;
wire n_16500;
wire n_16501;
wire n_16502;
wire n_16503;
wire n_16504;
wire n_16505;
wire n_16506;
wire n_16507;
wire n_16508;
wire n_16509;
wire n_16510;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16514;
wire n_16515;
wire n_16516;
wire n_16517;
wire n_16518;
wire n_16519;
wire n_16520;
wire n_16521;
wire n_16522;
wire n_16523;
wire n_16524;
wire n_16525;
wire n_16526;
wire n_16527;
wire n_16528;
wire n_16529;
wire n_16530;
wire n_16531;
wire n_16532;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16545;
wire n_16546;
wire n_16547;
wire n_16548;
wire n_16549;
wire n_16550;
wire n_16551;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_16555;
wire n_16556;
wire n_16557;
wire n_16558;
wire n_16559;
wire n_16560;
wire n_16561;
wire n_16562;
wire n_16563;
wire n_16564;
wire n_16565;
wire n_16566;
wire n_16567;
wire n_16568;
wire n_16569;
wire n_16570;
wire n_16571;
wire n_16572;
wire n_16573;
wire n_16574;
wire n_16575;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_16580;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_16590;
wire n_16591;
wire n_16592;
wire n_16593;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16598;
wire n_16599;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16604;
wire n_16605;
wire n_16606;
wire n_16607;
wire n_16608;
wire n_16609;
wire n_16610;
wire n_16611;
wire n_16612;
wire n_16613;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_16618;
wire n_16619;
wire n_16620;
wire n_16621;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire n_16626;
wire n_16627;
wire n_16628;
wire n_16629;
wire n_16630;
wire n_16631;
wire n_16632;
wire n_16633;
wire n_16634;
wire n_16635;
wire n_16636;
wire n_16637;
wire n_16638;
wire n_16639;
wire n_16640;
wire n_16641;
wire n_16642;
wire n_16643;
wire n_16644;
wire n_16645;
wire n_16646;
wire n_16647;
wire n_16648;
wire n_16649;
wire n_16650;
wire n_16651;
wire n_16652;
wire n_16653;
wire n_16654;
wire n_16655;
wire n_16656;
wire n_16657;
wire n_16658;
wire n_16659;
wire n_16660;
wire n_16661;
wire n_16662;
wire n_16663;
wire n_16664;
wire n_16665;
wire n_16666;
wire n_16667;
wire n_16668;
wire n_16669;
wire n_16670;
wire n_16671;
wire n_16672;
wire n_16673;
wire n_16674;
wire n_16675;
wire n_16676;
wire n_16677;
wire n_16678;
wire n_16679;
wire n_16680;
wire n_16681;
wire n_16682;
wire n_16683;
wire n_16684;
wire n_16685;
wire n_16686;
wire n_16687;
wire n_16688;
wire n_16689;
wire n_16690;
wire n_16691;
wire n_16692;
wire n_16693;
wire n_16694;
wire n_16695;
wire n_16696;
wire n_16697;
wire n_16698;
wire n_16699;
wire n_16700;
wire n_16701;
wire n_16702;
wire n_16703;
wire n_16704;
wire n_16705;
wire n_16706;
wire n_16707;
wire n_16708;
wire n_16709;
wire n_16710;
wire n_16711;
wire n_16712;
wire n_16713;
wire n_16714;
wire n_16715;
wire n_16716;
wire n_16717;
wire n_16718;
wire n_16719;
wire n_16720;
wire n_16721;
wire n_16722;
wire n_16723;
wire n_16724;
wire n_16725;
wire n_16726;
wire n_16727;
wire n_16728;
wire n_16729;
wire n_16730;
wire n_16731;
wire n_16732;
wire n_16733;
wire n_16734;
wire n_16735;
wire n_16736;
wire n_16737;
wire n_16738;
wire n_16739;
wire n_16740;
wire n_16741;
wire n_16742;
wire n_16743;
wire n_16744;
wire n_16745;
wire n_16746;
wire n_16747;
wire n_16748;
wire n_16749;
wire n_16750;
wire n_16751;
wire n_16752;
wire n_16753;
wire n_16754;
wire n_16755;
wire n_16756;
wire n_16757;
wire n_16758;
wire n_16759;
wire n_16760;
wire n_16761;
wire n_16762;
wire n_16763;
wire n_16764;
wire n_16765;
wire n_16766;
wire n_16767;
wire n_16768;
wire n_16769;
wire n_16770;
wire n_16771;
wire n_16772;
wire n_16773;
wire n_16774;
wire n_16775;
wire n_16776;
wire n_16777;
wire n_16778;
wire n_16779;
wire n_16780;
wire n_16781;
wire n_16782;
wire n_16783;
wire n_16784;
wire n_16785;
wire n_16786;
wire n_16787;
wire n_16788;
wire n_16789;
wire n_16790;
wire n_16791;
wire n_16792;
wire n_16793;
wire n_16794;
wire n_16795;
wire n_16796;
wire n_16797;
wire n_16798;
wire n_16799;
wire n_16800;
wire n_16801;
wire n_16802;
wire n_16803;
wire n_16804;
wire n_16805;
wire n_16806;
wire n_16807;
wire n_16808;
wire n_16809;
wire n_16810;
wire n_16811;
wire n_16812;
wire n_16813;
wire n_16814;
wire n_16815;
wire n_16816;
wire n_16817;
wire n_16818;
wire n_16819;
wire n_16820;
wire n_16821;
wire n_16822;
wire n_16823;
wire n_16824;
wire n_16825;
wire n_16826;
wire n_16827;
wire n_16828;
wire n_16829;
wire n_16830;
wire n_16831;
wire n_16832;
wire n_16833;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16846;
wire n_16847;
wire n_16848;
wire n_16849;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_16856;
wire n_16857;
wire n_16858;
wire n_16859;
wire n_16860;
wire n_16861;
wire n_16862;
wire n_16863;
wire n_16864;
wire n_16865;
wire n_16866;
wire n_16867;
wire n_16868;
wire n_16869;
wire n_16870;
wire n_16871;
wire n_16872;
wire n_16873;
wire n_16874;
wire n_16875;
wire n_16876;
wire n_16877;
wire n_16878;
wire n_16879;
wire n_16880;
wire n_16881;
wire n_16882;
wire n_16883;
wire n_16884;
wire n_16885;
wire n_16886;
wire n_16887;
wire n_16888;
wire n_16889;
wire n_16890;
wire n_16891;
wire n_16892;
wire n_16893;
wire n_16894;
wire n_16895;
wire n_16896;
wire n_16897;
wire n_16898;
wire n_16899;
wire n_16900;
wire n_16901;
wire n_16902;
wire n_16903;
wire n_16904;
wire n_16905;
wire n_16906;
wire n_16907;
wire n_16908;
wire n_16909;
wire n_16910;
wire n_16911;
wire n_16912;
wire n_16913;
wire n_16914;
wire n_16915;
wire n_16916;
wire n_16917;
wire n_16918;
wire n_16919;
wire n_16920;
wire n_16921;
wire n_16922;
wire n_16923;
wire n_16924;
wire n_16925;
wire n_16926;
wire n_16927;
wire n_16928;
wire n_16929;
wire n_16930;
wire n_16931;
wire n_16932;
wire n_16933;
wire n_16934;
wire n_16935;
wire n_16936;
wire n_16937;
wire n_16938;
wire n_16939;
wire n_16940;
wire n_16941;
wire n_16942;
wire n_16943;
wire n_16944;
wire n_16945;
wire n_16946;
wire n_16947;
wire n_16948;
wire n_16949;
wire n_16950;
wire n_16951;
wire n_16952;
wire n_16953;
wire n_16954;
wire n_16955;
wire n_16956;
wire n_16957;
wire n_16958;
wire n_16959;
wire n_16960;
wire n_16961;
wire n_16962;
wire n_16963;
wire n_16964;
wire n_16965;
wire n_16966;
wire n_16967;
wire n_16968;
wire n_16969;
wire n_16970;
wire n_16971;
wire n_16972;
wire n_16973;
wire n_16974;
wire n_16975;
wire n_16976;
wire n_16977;
wire n_16978;
wire n_16979;
wire n_16980;
wire n_16981;
wire n_16982;
wire n_16983;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_16988;
wire n_16989;
wire n_16990;
wire n_16991;
wire n_16992;
wire n_16993;
wire n_16994;
wire n_16995;
wire n_16996;
wire n_16997;
wire n_16998;
wire n_16999;
wire n_17000;
wire n_17001;
wire n_17002;
wire n_17003;
wire n_17004;
wire n_17005;
wire n_17006;
wire n_17007;
wire n_17008;
wire n_17009;
wire n_17010;
wire n_17011;
wire n_17012;
wire n_17013;
wire n_17014;
wire n_17015;
wire n_17016;
wire n_17017;
wire n_17018;
wire n_17019;
wire n_17020;
wire n_17021;
wire n_17022;
wire n_17023;
wire n_17024;
wire n_17025;
wire n_17026;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17033;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17037;
wire n_17038;
wire n_17039;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17047;
wire n_17048;
wire n_17049;
wire n_17050;
wire n_17051;
wire n_17052;
wire n_17053;
wire n_17054;
wire n_17055;
wire n_17056;
wire n_17057;
wire n_17058;
wire n_17059;
wire n_17060;
wire n_17061;
wire n_17062;
wire n_17063;
wire n_17064;
wire n_17065;
wire n_17066;
wire n_17067;
wire n_17068;
wire n_17069;
wire n_17070;
wire n_17071;
wire n_17072;
wire n_17073;
wire n_17074;
wire n_17075;
wire n_17076;
wire n_17077;
wire n_17078;
wire n_17079;
wire n_17080;
wire n_17081;
wire n_17082;
wire n_17083;
wire n_17084;
wire n_17085;
wire n_17086;
wire n_17087;
wire n_17088;
wire n_17089;
wire n_17090;
wire n_17091;
wire n_17092;
wire n_17093;
wire n_17094;
wire n_17095;
wire n_17096;
wire n_17097;
wire n_17098;
wire n_17099;
wire n_17100;
wire n_17101;
wire n_17102;
wire n_17103;
wire n_17104;
wire n_17105;
wire n_17106;
wire n_17107;
wire n_17108;
wire n_17109;
wire n_17110;
wire n_17111;
wire n_17112;
wire n_17113;
wire n_17114;
wire n_17115;
wire n_17116;
wire n_17117;
wire n_17118;
wire n_17119;
wire n_17120;
wire n_17121;
wire n_17122;
wire n_17123;
wire n_17124;
wire n_17125;
wire n_17126;
wire n_17127;
wire n_17128;
wire n_17129;
wire n_17130;
wire n_17131;
wire n_17132;
wire n_17133;
wire n_17134;
wire n_17135;
wire n_17136;
wire n_17137;
wire n_17138;
wire n_17139;
wire n_17140;
wire n_17141;
wire n_17142;
wire n_17143;
wire n_17144;
wire n_17145;
wire n_17146;
wire n_17147;
wire n_17148;
wire n_17149;
wire n_17150;
wire n_17151;
wire n_17152;
wire n_17153;
wire n_17154;
wire n_17155;
wire n_17156;
wire n_17157;
wire n_17158;
wire n_17159;
wire n_17160;
wire n_17161;
wire n_17162;
wire n_17163;
wire n_17164;
wire n_17165;
wire n_17166;
wire n_17167;
wire n_17168;
wire n_17169;
wire n_17170;
wire n_17171;
wire n_17172;
wire n_17173;
wire n_17174;
wire n_17175;
wire n_17176;
wire n_17177;
wire n_17178;
wire n_17179;
wire n_17180;
wire n_17181;
wire n_17182;
wire n_17183;
wire n_17184;
wire n_17185;
wire n_17186;
wire n_17187;
wire n_17188;
wire n_17189;
wire n_17190;
wire n_17191;
wire n_17192;
wire n_17193;
wire n_17194;
wire n_17195;
wire n_17196;
wire n_17197;
wire n_17198;
wire n_17199;
wire n_17200;
wire n_17201;
wire n_17202;
wire n_17203;
wire n_17204;
wire n_17205;
wire n_17206;
wire n_17207;
wire n_17208;
wire n_17209;
wire n_17210;
wire n_17211;
wire n_17212;
wire n_17213;
wire n_17214;
wire n_17215;
wire n_17216;
wire n_17217;
wire n_17218;
wire n_17219;
wire n_17220;
wire n_17221;
wire n_17222;
wire n_17223;
wire n_17224;
wire n_17225;
wire n_17226;
wire n_17227;
wire n_17228;
wire n_17229;
wire n_17230;
wire n_17231;
wire n_17232;
wire n_17233;
wire n_17234;
wire n_17235;
wire n_17236;
wire n_17237;
wire n_17238;
wire n_17239;
wire n_17240;
wire n_17241;
wire n_17242;
wire n_17243;
wire n_17244;
wire n_17245;
wire n_17246;
wire n_17247;
wire n_17248;
wire n_17249;
wire n_17250;
wire n_17251;
wire n_17252;
wire n_17253;
wire n_17254;
wire n_17255;
wire n_17256;
wire n_17257;
wire n_17258;
wire n_17259;
wire n_17260;
wire n_17261;
wire n_17262;
wire n_17263;
wire n_17264;
wire n_17265;
wire n_17266;
wire n_17267;
wire n_17268;
wire n_17269;
wire n_17270;
wire n_17271;
wire n_17272;
wire n_17273;
wire n_17274;
wire n_17275;
wire n_17276;
wire n_17277;
wire n_17278;
wire n_17279;
wire n_17280;
wire n_17281;
wire n_17282;
wire n_17283;
wire n_17284;
wire n_17285;
wire n_17286;
wire n_17287;
wire n_17288;
wire n_17289;
wire n_17290;
wire n_17291;
wire n_17292;
wire n_17293;
wire n_17294;
wire n_17295;
wire n_17296;
wire n_17297;
wire n_17298;
wire n_17299;
wire n_17300;
wire n_17301;
wire n_17302;
wire n_17303;
wire n_17304;
wire n_17305;
wire n_17306;
wire n_17307;
wire n_17308;
wire n_17309;
wire n_17310;
wire n_17311;
wire n_17312;
wire n_17313;
wire n_17314;
wire n_17315;
wire n_17316;
wire n_17317;
wire n_17318;
wire n_17319;
wire n_17320;
wire n_17321;
wire n_17322;
wire n_17323;
wire n_17324;
wire n_17325;
wire n_17326;
wire n_17327;
wire n_17328;
wire n_17329;
wire n_17330;
wire n_17331;
wire n_17332;
wire n_17333;
wire n_17334;
wire n_17335;
wire n_17336;
wire n_17337;
wire n_17338;
wire n_17339;
wire n_17340;
wire n_17341;
wire n_17342;
wire n_17343;
wire n_17344;
wire n_17345;
wire n_17346;
wire n_17347;
wire n_17348;
wire n_17349;
wire n_17350;
wire n_17351;
wire n_17352;
wire n_17353;
wire n_17354;
wire n_17355;
wire n_17356;
wire n_17357;
wire n_17358;
wire n_17359;
wire n_17360;
wire n_17361;
wire n_17362;
wire n_17363;
wire n_17364;
wire n_17365;
wire n_17366;
wire n_17367;
wire n_17368;
wire n_17369;
wire n_17370;
wire n_17371;
wire n_17372;
wire n_17373;
wire n_17374;
wire n_17375;
wire n_17376;
wire n_17377;
wire n_17378;
wire n_17379;
wire n_17380;
wire n_17381;
wire n_17382;
wire n_17383;
wire n_17384;
wire n_17385;
wire n_17386;
wire n_17387;
wire n_17388;
wire n_17389;
wire n_17390;
wire n_17391;
wire n_17392;
wire n_17393;
wire n_17394;
wire n_17395;
wire n_17396;
wire n_17397;
wire n_17398;
wire n_17399;
wire n_17400;
wire n_17401;
wire n_17402;
wire n_17403;
wire n_17404;
wire n_17405;
wire n_17406;
wire n_17407;
wire n_17408;
wire n_17409;
wire n_17410;
wire n_17411;
wire n_17412;
wire n_17413;
wire n_17414;
wire n_17415;
wire n_17416;
wire n_17417;
wire n_17418;
wire n_17419;
wire n_17420;
wire n_17421;
wire n_17422;
wire n_17423;
wire n_17424;
wire n_17425;
wire n_17426;
wire n_17427;
wire n_17428;
wire n_17429;
wire n_17430;
wire n_17431;
wire n_17432;
wire n_17433;
wire n_17434;
wire n_17435;
wire n_17436;
wire n_17437;
wire n_17438;
wire n_17439;
wire n_17440;
wire n_17441;
wire n_17442;
wire n_17443;
wire n_17444;
wire n_17445;
wire n_17446;
wire n_17447;
wire n_17448;
wire n_17449;
wire n_17450;
wire n_17451;
wire n_17452;
wire n_17453;
wire n_17454;
wire n_17455;
wire n_17456;
wire n_17457;
wire n_17458;
wire n_17459;
wire n_17460;
wire n_17461;
wire n_17462;
wire n_17463;
wire n_17464;
wire n_17465;
wire n_17466;
wire n_17467;
wire n_17468;
wire n_17469;
wire n_17470;
wire n_17471;
wire n_17472;
wire n_17473;
wire n_17474;
wire n_17475;
wire n_17476;
wire n_17477;
wire n_17478;
wire n_17479;
wire n_17480;
wire n_17481;
wire n_17482;
wire n_17483;
wire n_17484;
wire n_17485;
wire n_17486;
wire n_17487;
wire n_17488;
wire n_17489;
wire n_17490;
wire n_17491;
wire n_17492;
wire n_17493;
wire n_17494;
wire n_17495;
wire n_17496;
wire n_17497;
wire n_17498;
wire n_17499;
wire n_17500;
wire n_17501;
wire n_17502;
wire n_17503;
wire n_17504;
wire n_17505;
wire n_17506;
wire n_17507;
wire n_17508;
wire n_17509;
wire n_17510;
wire n_17511;
wire n_17512;
wire n_17513;
wire n_17514;
wire n_17515;
wire n_17516;
wire n_17517;
wire n_17518;
wire n_17519;
wire n_17520;
wire n_17521;
wire n_17522;
wire n_17523;
wire n_17524;
wire n_17525;
wire n_17526;
wire n_17527;
wire n_17528;
wire n_17529;
wire n_17530;
wire n_17531;
wire n_17532;
wire n_17533;
wire n_17534;
wire n_17535;
wire n_17536;
wire n_17537;
wire n_17538;
wire n_17539;
wire n_17540;
wire n_17541;
wire n_17542;
wire n_17543;
wire n_17544;
wire n_17545;
wire n_17546;
wire n_17547;
wire n_17548;
wire n_17549;
wire n_17550;
wire n_17551;
wire n_17552;
wire n_17553;
wire n_17554;
wire n_17555;
wire n_17556;
wire n_17557;
wire n_17558;
wire n_17559;
wire n_17560;
wire n_17561;
wire n_17562;
wire n_17563;
wire n_17564;
wire n_17565;
wire n_17566;
wire n_17567;
wire n_17568;
wire n_17569;
wire n_17570;
wire n_17571;
wire n_17572;
wire n_17573;
wire n_17574;
wire n_17575;
wire n_17576;
wire n_17577;
wire n_17578;
wire n_17579;
wire n_17580;
wire n_17581;
wire n_17582;
wire n_17583;
wire n_17584;
wire n_17585;
wire n_17586;
wire n_17587;
wire n_17588;
wire n_17589;
wire n_17590;
wire n_17591;
wire n_17592;
wire n_17593;
wire n_17594;
wire n_17595;
wire n_17596;
wire n_17597;
wire n_17598;
wire n_17599;
wire n_17600;
wire n_17601;
wire n_17602;
wire n_17603;
wire n_17604;
wire n_17605;
wire n_17606;
wire n_17607;
wire n_17608;
wire n_17609;
wire n_17610;
wire n_17611;
wire n_17612;
wire n_17613;
wire n_17614;
wire n_17615;
wire n_17616;
wire n_17617;
wire n_17618;
wire n_17619;
wire n_17620;
wire n_17621;
wire n_17622;
wire n_17623;
wire n_17624;
wire n_17625;
wire n_17626;
wire n_17627;
wire n_17628;
wire n_17629;
wire n_17630;
wire n_17631;
wire n_17632;
wire n_17633;
wire n_17634;
wire n_17635;
wire n_17636;
wire n_17637;
wire n_17638;
wire n_17639;
wire n_17640;
wire n_17641;
wire n_17642;
wire n_17643;
wire n_17644;
wire n_17645;
wire n_17646;
wire n_17647;
wire n_17648;
wire n_17649;
wire n_17650;
wire n_17651;
wire n_17652;
wire n_17653;
wire n_17654;
wire n_17655;
wire n_17656;
wire n_17657;
wire n_17658;
wire n_17659;
wire n_17660;
wire n_17661;
wire n_17662;
wire n_17663;
wire n_17664;
wire n_17665;
wire n_17666;
wire n_17667;
wire n_17668;
wire n_17669;
wire n_17670;
wire n_17671;
wire n_17672;
wire n_17673;
wire n_17674;
wire n_17675;
wire n_17676;
wire n_17677;
wire n_17678;
wire n_17679;
wire n_17680;
wire n_17681;
wire n_17682;
wire n_17683;
wire n_17684;
wire n_17685;
wire n_17686;
wire n_17687;
wire n_17688;
wire n_17689;
wire n_17690;
wire n_17691;
wire n_17692;
wire n_17693;
wire n_17694;
wire n_17695;
wire n_17696;
wire n_17697;
wire n_17698;
wire n_17699;
wire n_17700;
wire n_17701;
wire n_17702;
wire n_17703;
wire n_17704;
wire n_17705;
wire n_17706;
wire n_17707;
wire n_17708;
wire n_17709;
wire n_17710;
wire n_17711;
wire n_17712;
wire n_17713;
wire n_17714;
wire n_17715;
wire n_17716;
wire n_17717;
wire n_17718;
wire n_17719;
wire n_17720;
wire n_17721;
wire n_17722;
wire n_17723;
wire n_17724;
wire n_17725;
wire n_17726;
wire n_17727;
wire n_17728;
wire n_17729;
wire n_17730;
wire n_17731;
wire n_17732;
wire n_17733;
wire n_17734;
wire n_17735;
wire n_17736;
wire n_17737;
wire n_17738;
wire n_17739;
wire n_17740;
wire n_17741;
wire n_17742;
wire n_17743;
wire n_17744;
wire n_17745;
wire n_17746;
wire n_17747;
wire n_17748;
wire n_17749;
wire n_17750;
wire n_17751;
wire n_17752;
wire n_17753;
wire n_17754;
wire n_17755;
wire n_17756;
wire n_17757;
wire n_17758;
wire n_17759;
wire n_17760;
wire n_17761;
wire n_17762;
wire n_17763;
wire n_17764;
wire n_17765;
wire n_17766;
wire n_17767;
wire n_17768;
wire n_17769;
wire n_17770;
wire n_17771;
wire n_17772;
wire n_17773;
wire n_17774;
wire n_17775;
wire n_17776;
wire n_17777;
wire n_17778;
wire n_17779;
wire n_17780;
wire n_17781;
wire n_17782;
wire n_17783;
wire n_17784;
wire n_17785;
wire n_17786;
wire n_17787;
wire n_17788;
wire n_17789;
wire n_17790;
wire n_17791;
wire n_17792;
wire n_17793;
wire n_17794;
wire n_17795;
wire n_17796;
wire n_17797;
wire n_17798;
wire n_17799;
wire n_17800;
wire n_17801;
wire n_17802;
wire n_17803;
wire n_17804;
wire n_17805;
wire n_17806;
wire n_17807;
wire n_17808;
wire n_17809;
wire n_17810;
wire n_17811;
wire n_17812;
wire n_17813;
wire n_17814;
wire n_17815;
wire n_17816;
wire n_17817;
wire n_17818;
wire n_17819;
wire n_17820;
wire n_17821;
wire n_17822;
wire n_17823;
wire n_17824;
wire n_17825;
wire n_17826;
wire n_17827;
wire n_17828;
wire n_17829;
wire n_17830;
wire n_17831;
wire n_17832;
wire n_17833;
wire n_17834;
wire n_17835;
wire n_17836;
wire n_17837;
wire n_17838;
wire n_17839;
wire n_17840;
wire n_17841;
wire n_17842;
wire n_17843;
wire n_17844;
wire n_17845;
wire n_17846;
wire n_17847;
wire n_17848;
wire n_17849;
wire n_17850;
wire n_17851;
wire n_17852;
wire n_17853;
wire n_17854;
wire n_17855;
wire n_17856;
wire n_17857;
wire n_17858;
wire n_17859;
wire n_17860;
wire n_17861;
wire n_17862;
wire n_17863;
wire n_17864;
wire n_17865;
wire n_17866;
wire n_17867;
wire n_17868;
wire n_17869;
wire n_17870;
wire n_17871;
wire n_17872;
wire n_17873;
wire n_17874;
wire n_17875;
wire n_17876;
wire n_17877;
wire n_17878;
wire n_17879;
wire n_17880;
wire n_17881;
wire n_17882;
wire n_17883;
wire n_17884;
wire n_17885;
wire n_17886;
wire n_17887;
wire n_17888;
wire n_17889;
wire n_17890;
wire n_17891;
wire n_17892;
wire n_17893;
wire n_17894;
wire n_17895;
wire n_17896;
wire n_17897;
wire n_17898;
wire n_17899;
wire n_17900;
wire n_17901;
wire n_17902;
wire n_17903;
wire n_17904;
wire n_17905;
wire n_17906;
wire n_17907;
wire n_17908;
wire n_17909;
wire n_17910;
wire n_17911;
wire n_17912;
wire n_17913;
wire n_17914;
wire n_17915;
wire n_17916;
wire n_17917;
wire n_17918;
wire n_17919;
wire n_17920;
wire n_17921;
wire n_17922;
wire n_17923;
wire n_17924;
wire n_17925;
wire n_17926;
wire n_17927;
wire n_17928;
wire n_17929;
wire n_17930;
wire n_17931;
wire n_17932;
wire n_17933;
wire n_17934;
wire n_17935;
wire n_17936;
wire n_17937;
wire n_17938;
wire n_17939;
wire n_17940;
wire n_17941;
wire n_17942;
wire n_17943;
wire n_17944;
wire n_17945;
wire n_17946;
wire n_17947;
wire n_17948;
wire n_17949;
wire n_17950;
wire n_17951;
wire n_17952;
wire n_17953;
wire n_17954;
wire n_17955;
wire n_17956;
wire n_17957;
wire n_17958;
wire n_17959;
wire n_17960;
wire n_17961;
wire n_17962;
wire n_17963;
wire n_17964;
wire n_17965;
wire n_17966;
wire n_17967;
wire n_17968;
wire n_17969;
wire n_17970;
wire n_17971;
wire n_17972;
wire n_17973;
wire n_17974;
wire n_17975;
wire n_17976;
wire n_17977;
wire n_17978;
wire n_17979;
wire n_17980;
wire n_17981;
wire n_17982;
wire n_17983;
wire n_17984;
wire n_17985;
wire n_17986;
wire n_17987;
wire n_17988;
wire n_17989;
wire n_17990;
wire n_17991;
wire n_17992;
wire n_17993;
wire n_17994;
wire n_17995;
wire n_17996;
wire n_17997;
wire n_17998;
wire n_17999;
wire n_18000;
wire n_18001;
wire n_18002;
wire n_18003;
wire n_18004;
wire n_18005;
wire n_18006;
wire n_18007;
wire n_18008;
wire n_18009;
wire n_18010;
wire n_18011;
wire n_18012;
wire n_18013;
wire n_18014;
wire n_18015;
wire n_18016;
wire n_18017;
wire n_18018;
wire n_18019;
wire n_18020;
wire n_18021;
wire n_18022;
wire n_18023;
wire n_18024;
wire n_18025;
wire n_18026;
wire n_18027;
wire n_18028;
wire n_18029;
wire n_18030;
wire n_18031;
wire n_18032;
wire n_18033;
wire n_18034;
wire n_18035;
wire n_18036;
wire n_18037;
wire n_18038;
wire n_18039;
wire n_18040;
wire n_18041;
wire n_18042;
wire n_18043;
wire n_18044;
wire n_18045;
wire n_18046;
wire n_18047;
wire n_18048;
wire n_18049;
wire n_18050;
wire n_18051;
wire n_18052;
wire n_18053;
wire n_18054;
wire n_18055;
wire n_18056;
wire n_18057;
wire n_18058;
wire n_18059;
wire n_18060;
wire n_18061;
wire n_18062;
wire n_18063;
wire n_18064;
wire n_18065;
wire n_18066;
wire n_18067;
wire n_18068;
wire n_18069;
wire n_18070;
wire n_18071;
wire n_18072;
wire n_18073;
wire n_18074;
wire n_18075;
wire n_18076;
wire n_18077;
wire n_18078;
wire n_18079;
wire n_18080;
wire n_18081;
wire n_18082;
wire n_18083;
wire n_18084;
wire n_18085;
wire n_18086;
wire n_18087;
wire n_18088;
wire n_18089;
wire n_18090;
wire n_18091;
wire n_18092;
wire n_18093;
wire n_18094;
wire n_18095;
wire n_18096;
wire n_18097;
wire n_18098;
wire n_18099;
wire n_18100;
wire n_18101;
wire n_18102;
wire n_18103;
wire n_18104;
wire n_18105;
wire n_18106;
wire n_18107;
wire n_18108;
wire n_18109;
wire n_18110;
wire n_18111;
wire n_18112;
wire n_18113;
wire n_18114;
wire n_18115;
wire n_18116;
wire n_18117;
wire n_18118;
wire n_18119;
wire n_18120;
wire n_18121;
wire n_18122;
wire n_18123;
wire n_18124;
wire n_18125;
wire n_18126;
wire n_18127;
wire n_18128;
wire n_18129;
wire n_18130;
wire n_18131;
wire n_18132;
wire n_18133;
wire n_18134;
wire n_18135;
wire n_18136;
wire n_18137;
wire n_18138;
wire n_18139;
wire n_18140;
wire n_18141;
wire n_18142;
wire n_18143;
wire n_18144;
wire n_18145;
wire n_18146;
wire n_18147;
wire n_18148;
wire n_18149;
wire n_18150;
wire n_18151;
wire n_18152;
wire n_18153;
wire n_18154;
wire n_18155;
wire n_18156;
wire n_18157;
wire n_18158;
wire n_18159;
wire n_18160;
wire n_18161;
wire n_18162;
wire n_18163;
wire n_18164;
wire n_18165;
wire n_18166;
wire n_18167;
wire n_18168;
wire n_18169;
wire n_18170;
wire n_18171;
wire n_18172;
wire n_18173;
wire n_18174;
wire n_18175;
wire n_18176;
wire n_18177;
wire n_18178;
wire n_18179;
wire n_18180;
wire n_18181;
wire n_18182;
wire n_18183;
wire n_18184;
wire n_18185;
wire n_18186;
wire n_18187;
wire n_18188;
wire n_18189;
wire n_18190;
wire n_18191;
wire n_18192;
wire n_18193;
wire n_18194;
wire n_18195;
wire n_18196;
wire n_18197;
wire n_18198;
wire n_18199;
wire n_18200;
wire n_18201;
wire n_18202;
wire n_18203;
wire n_18204;
wire n_18205;
wire n_18206;
wire n_18207;
wire n_18208;
wire n_18209;
wire n_18210;
wire n_18211;
wire n_18212;
wire n_18213;
wire n_18214;
wire n_18215;
wire n_18216;
wire n_18217;
wire n_18218;
wire n_18219;
wire n_18220;
wire n_18221;
wire n_18222;
wire n_18223;
wire n_18224;
wire n_18225;
wire n_18226;
wire n_18227;
wire n_18228;
wire n_18229;
wire n_18230;
wire n_18231;
wire n_18232;
wire n_18233;
wire n_18234;
wire n_18235;
wire n_18236;
wire n_18237;
wire n_18238;
wire n_18239;
wire n_18240;
wire n_18241;
wire n_18242;
wire n_18243;
wire n_18244;
wire n_18245;
wire n_18246;
wire n_18247;
wire n_18248;
wire n_18249;
wire n_18250;
wire n_18251;
wire n_18252;
wire n_18253;
wire n_18254;
wire n_18255;
wire n_18256;
wire n_18257;
wire n_18258;
wire n_18259;
wire n_18260;
wire n_18261;
wire n_18262;
wire n_18263;
wire n_18264;
wire n_18265;
wire n_18266;
wire n_18267;
wire n_18268;
wire n_18269;
wire n_18270;
wire n_18271;
wire n_18272;
wire n_18273;
wire n_18274;
wire n_18275;
wire n_18276;
wire n_18277;
wire n_18278;
wire n_18279;
wire n_18280;
wire n_18281;
wire n_18282;
wire n_18283;
wire n_18284;
wire n_18285;
wire n_18286;
wire n_18287;
wire n_18288;
wire n_18289;
wire n_18290;
wire n_18291;
wire n_18292;
wire n_18293;
wire n_18294;
wire n_18295;
wire n_18296;
wire n_18297;
wire n_18298;
wire n_18299;
wire n_18300;
wire n_18301;
wire n_18302;
wire n_18303;
wire n_18304;
wire n_18305;
wire n_18306;
wire n_18307;
wire n_18308;
wire n_18309;
wire n_18310;
wire n_18311;
wire n_18312;
wire n_18313;
wire n_18314;
wire n_18315;
wire n_18316;
wire n_18317;
wire n_18318;
wire n_18319;
wire n_18320;
wire n_18321;
wire n_18322;
wire n_18323;
wire n_18324;
wire n_18325;
wire n_18326;
wire n_18327;
wire n_18328;
wire n_18329;
wire n_18330;
wire n_18331;
wire n_18332;
wire n_18333;
wire n_18334;
wire n_18335;
wire n_18336;
wire n_18337;
wire n_18338;
wire n_18339;
wire n_18340;
wire n_18341;
wire n_18342;
wire n_18343;
wire n_18344;
wire n_18345;
wire n_18346;
wire n_18347;
wire n_18348;
wire n_18349;
wire n_18350;
wire n_18351;
wire n_18352;
wire n_18353;
wire n_18354;
wire n_18355;
wire n_18356;
wire n_18357;
wire n_18358;
wire n_18359;
wire n_18360;
wire n_18361;
wire n_18362;
wire n_18363;
wire n_18364;
wire n_18365;
wire n_18366;
wire n_18367;
wire n_18368;
wire n_18369;
wire n_18370;
wire n_18371;
wire n_18372;
wire n_18373;
wire n_18374;
wire n_18375;
wire n_18376;
wire n_18377;
wire n_18378;
wire n_18379;
wire n_18380;
wire n_18381;
wire n_18382;
wire n_18383;
wire n_18384;
wire n_18385;
wire n_18386;
wire n_18387;
wire n_18388;
wire n_18389;
wire n_18390;
wire n_18391;
wire n_18392;
wire n_18393;
wire n_18394;
wire n_18395;
wire n_18396;
wire n_18397;
wire n_18398;
wire n_18399;
wire n_18400;
wire n_18401;
wire n_18402;
wire n_18403;
wire n_18404;
wire n_18405;
wire n_18406;
wire n_18407;
wire n_18408;
wire n_18409;
wire n_18410;
wire n_18411;
wire n_18412;
wire n_18413;
wire n_18414;
wire n_18415;
wire n_18416;
wire n_18417;
wire n_18418;
wire n_18419;
wire n_18420;
wire n_18421;
wire n_18422;
wire n_18423;
wire n_18424;
wire n_18425;
wire n_18426;
wire n_18427;
wire n_18428;
wire n_18429;
wire n_18430;
wire n_18431;
wire n_18432;
wire n_18433;
wire n_18434;
wire n_18435;
wire n_18436;
wire n_18437;
wire n_18438;
wire n_18439;
wire n_18440;
wire n_18441;
wire n_18442;
wire n_18443;
wire n_18444;
wire n_18445;
wire n_18446;
wire n_18447;
wire n_18448;
wire n_18449;
wire n_18450;
wire n_18451;
wire n_18452;
wire n_18453;
wire n_18454;
wire n_18455;
wire n_18456;
wire n_18457;
wire n_18458;
wire n_18459;
wire n_18460;
wire n_18461;
wire n_18462;
wire n_18463;
wire n_18464;
wire n_18465;
wire n_18466;
wire n_18467;
wire n_18468;
wire n_18469;
wire n_18470;
wire n_18471;
wire n_18472;
wire n_18473;
wire n_18474;
wire n_18475;
wire n_18476;
wire n_18477;
wire n_18478;
wire n_18479;
wire n_18480;
wire n_18481;
wire n_18482;
wire n_18483;
wire n_18484;
wire n_18485;
wire n_18486;
wire n_18487;
wire n_18488;
wire n_18489;
wire n_18490;
wire n_18491;
wire n_18492;
wire n_18493;
wire n_18494;
wire n_18495;
wire n_18496;
wire n_18497;
wire n_18498;
wire n_18499;
wire n_18500;
wire n_18501;
wire n_18502;
wire n_18503;
wire n_18504;
wire n_18505;
wire n_18506;
wire n_18507;
wire n_18508;
wire n_18509;
wire n_18510;
wire n_18511;
wire n_18512;
wire n_18513;
wire n_18514;
wire n_18515;
wire n_18516;
wire n_18517;
wire n_18518;
wire n_18519;
wire n_18520;
wire n_18521;
wire n_18522;
wire n_18523;
wire n_18524;
wire n_18525;
wire n_18526;
wire n_18527;
wire n_18528;
wire n_18529;
wire n_18530;
wire n_18531;
wire n_18532;
wire n_18533;
wire n_18534;
wire n_18535;
wire n_18536;
wire n_18537;
wire n_18538;
wire n_18539;
wire n_18540;
wire n_18541;
wire n_18542;
wire n_18543;
wire n_18544;
wire n_18545;
wire n_18546;
wire n_18547;
wire n_18548;
wire n_18549;
wire n_18550;
wire n_18551;
wire n_18552;
wire n_18553;
wire n_18554;
wire n_18555;
wire n_18556;
wire n_18557;
wire n_18558;
wire n_18559;
wire n_18560;
wire n_18561;
wire n_18562;
wire n_18563;
wire n_18564;
wire n_18565;
wire n_18566;
wire n_18567;
wire n_18568;
wire n_18569;
wire n_18570;
wire n_18571;
wire n_18572;
wire n_18573;
wire n_18574;
wire n_18575;
wire n_18576;
wire n_18577;
wire n_18578;
wire n_18579;
wire n_18580;
wire n_18581;
wire n_18582;
wire n_18583;
wire n_18584;
wire n_18585;
wire n_18586;
wire n_18587;
wire n_18588;
wire n_18589;
wire n_18590;
wire n_18591;
wire n_18592;
wire n_18593;
wire n_18594;
wire n_18595;
wire n_18596;
wire n_18597;
wire n_18598;
wire n_18599;
wire n_18600;
wire n_18601;
wire n_18602;
wire n_18603;
wire n_18604;
wire n_18605;
wire n_18606;
wire n_18607;
wire n_18608;
wire n_18609;
wire n_18610;
wire n_18611;
wire n_18612;
wire n_18613;
wire n_18614;
wire n_18615;
wire n_18616;
wire n_18617;
wire n_18618;
wire n_18619;
wire n_18620;
wire n_18621;
wire n_18622;
wire n_18623;
wire n_18624;
wire n_18625;
wire n_18626;
wire n_18627;
wire n_18628;
wire n_18629;
wire n_18630;
wire n_18631;
wire n_18632;
wire n_18633;
wire n_18634;
wire n_18635;
wire n_18636;
wire n_18637;
wire n_18638;
wire n_18639;
wire n_18640;
wire n_18641;
wire n_18642;
wire n_18643;
wire n_18644;
wire n_18645;
wire n_18646;
wire n_18647;
wire n_18648;
wire n_18649;
wire n_18650;
wire n_18651;
wire n_18652;
wire n_18653;
wire n_18654;
wire n_18655;
wire n_18656;
wire n_18657;
wire n_18658;
wire n_18659;
wire n_18660;
wire n_18661;
wire n_18662;
wire n_18663;
wire n_18664;
wire n_18665;
wire n_18666;
wire n_18667;
wire n_18668;
wire n_18669;
wire n_18670;
wire n_18671;
wire n_18672;
wire n_18673;
wire n_18674;
wire n_18675;
wire n_18676;
wire n_18677;
wire n_18678;
wire n_18679;
wire n_18680;
wire n_18681;
wire n_18682;
wire n_18683;
wire n_18684;
wire n_18685;
wire n_18686;
wire n_18687;
wire n_18688;
wire n_18689;
wire n_18690;
wire n_18691;
wire n_18692;
wire n_18693;
wire n_18694;
wire n_18695;
wire n_18696;
wire n_18697;
wire n_18698;
wire n_18699;
wire n_18700;
wire n_18701;
wire n_18702;
wire n_18703;
wire n_18704;
wire n_18705;
wire n_18706;
wire n_18707;
wire n_18708;
wire n_18709;
wire n_18710;
wire n_18711;
wire n_18712;
wire n_18713;
wire n_18714;
wire n_18715;
wire n_18716;
wire n_18717;
wire n_18718;
wire n_18719;
wire n_18720;
wire n_18721;
wire n_18722;
wire n_18723;
wire n_18724;
wire n_18725;
wire n_18726;
wire n_18727;
wire n_18728;
wire n_18729;
wire n_18730;
wire n_18731;
wire n_18732;
wire n_18733;
wire n_18734;
wire n_18735;
wire n_18736;
wire n_18737;
wire n_18738;
wire n_18739;
wire n_18740;
wire n_18741;
wire n_18742;
wire n_18743;
wire n_18744;
wire n_18745;
wire n_18746;
wire n_18747;
wire n_18748;
wire n_18749;
wire n_18750;
wire n_18751;
wire n_18752;
wire n_18753;
wire n_18754;
wire n_18755;
wire n_18756;
wire n_18757;
wire n_18758;
wire n_18759;
wire n_18760;
wire n_18761;
wire n_18762;
wire n_18763;
wire n_18764;
wire n_18765;
wire n_18766;
wire n_18767;
wire n_18768;
wire n_18769;
wire n_18770;
wire n_18771;
wire n_18772;
wire n_18773;
wire n_18774;
wire n_18775;
wire n_18776;
wire n_18777;
wire n_18778;
wire n_18779;
wire n_18780;
wire n_18781;
wire n_18782;
wire n_18783;
wire n_18784;
wire n_18785;
wire n_18786;
wire n_18787;
wire n_18788;
wire n_18789;
wire n_18790;
wire n_18791;
wire n_18792;
wire n_18793;
wire n_18794;
wire n_18795;
wire n_18796;
wire n_18797;
wire n_18798;
wire n_18799;
wire n_18800;
wire n_18801;
wire n_18802;
wire n_18803;
wire n_18804;
wire n_18805;
wire n_18806;
wire n_18807;
wire n_18808;
wire n_18809;
wire n_18810;
wire n_18811;
wire n_18812;
wire n_18813;
wire n_18814;
wire n_18815;
wire n_18816;
wire n_18817;
wire n_18818;
wire n_18819;
wire n_18820;
wire n_18821;
wire n_18822;
wire n_18823;
wire n_18824;
wire n_18825;
wire n_18826;
wire n_18827;
wire n_18828;
wire n_18829;
wire n_18830;
wire n_18831;
wire n_18832;
wire n_18833;
wire n_18834;
wire n_18835;
wire n_18836;
wire n_18837;
wire n_18838;
wire n_18839;
wire n_18840;
wire n_18841;
wire n_18842;
wire n_18843;
wire n_18844;
wire n_18845;
wire n_18846;
wire n_18847;
wire n_18848;
wire n_18849;
wire n_18850;
wire n_18851;
wire n_18852;
wire n_18853;
wire n_18854;
wire n_18855;
wire n_18856;
wire n_18857;
wire n_18858;
wire n_18859;
wire n_18860;
wire n_18861;
wire n_18862;
wire n_18863;
wire n_18864;
wire n_18865;
wire n_18866;
wire n_18867;
wire n_18868;
wire n_18869;
wire n_18870;
wire n_18871;
wire n_18872;
wire n_18873;
wire n_18874;
wire n_18875;
wire n_18876;
wire n_18877;
wire n_18878;
wire n_18879;
wire n_18880;
wire n_18881;
wire n_18882;
wire n_18883;
wire n_18884;
wire n_18885;
wire n_18886;
wire n_18887;
wire n_18888;
wire n_18889;
wire n_18890;
wire n_18891;
wire n_18892;
wire n_18893;
wire n_18894;
wire n_18895;
wire n_18896;
wire n_18897;
wire n_18898;
wire n_18899;
wire n_18900;
wire n_18901;
wire n_18902;
wire n_18903;
wire n_18904;
wire n_18905;
wire n_18906;
wire n_18907;
wire n_18908;
wire n_18909;
wire n_18910;
wire n_18911;
wire n_18912;
wire n_18913;
wire n_18914;
wire n_18915;
wire n_18916;
wire n_18917;
wire n_18918;
wire n_18919;
wire n_18920;
wire n_18921;
wire n_18922;
wire n_18923;
wire n_18924;
wire n_18925;
wire n_18926;
wire n_18927;
wire n_18928;
wire n_18929;
wire n_18930;
wire n_18931;
wire n_18932;
wire n_18933;
wire n_18934;
wire n_18935;
wire n_18936;
wire n_18937;
wire n_18938;
wire n_18939;
wire n_18940;
wire n_18941;
wire n_18942;
wire n_18943;
wire n_18944;
wire n_18945;
wire n_18946;
wire n_18947;
wire n_18948;
wire n_18949;
wire n_18950;
wire n_18951;
wire n_18952;
wire n_18953;
wire n_18954;
wire n_18955;
wire n_18956;
wire n_18957;
wire n_18958;
wire n_18959;
wire n_18960;
wire n_18961;
wire n_18962;
wire n_18963;
wire n_18964;
wire n_18965;
wire n_18966;
wire n_18967;
wire n_18968;
wire n_18969;
wire n_18970;
wire n_18971;
wire n_18972;
wire n_18973;
wire n_18974;
wire n_18975;
wire n_18976;
wire n_18977;
wire n_18978;
wire n_18979;
wire n_18980;
wire n_18981;
wire n_18982;
wire n_18983;
wire n_18984;
wire n_18985;
wire n_18986;
wire n_18987;
wire n_18988;
wire n_18989;
wire n_18990;
wire n_18991;
wire n_18992;
wire n_18993;
wire n_18994;
wire n_18995;
wire n_18996;
wire n_18997;
wire n_18998;
wire n_18999;
wire n_19000;
wire n_19001;
wire n_19002;
wire n_19003;
wire n_19004;
wire n_19005;
wire n_19006;
wire n_19007;
wire n_19008;
wire n_19009;
wire n_19010;
wire n_19011;
wire n_19012;
wire n_19013;
wire n_19014;
wire n_19015;
wire n_19016;
wire n_19017;
wire n_19018;
wire n_19019;
wire n_19020;
wire n_19021;
wire n_19022;
wire n_19023;
wire n_19024;
wire n_19025;
wire n_19026;
wire n_19027;
wire n_19028;
wire n_19029;
wire n_19030;
wire n_19031;
wire n_19032;
wire n_19033;
wire n_19034;
wire n_19035;
wire n_19036;
wire n_19037;
wire n_19038;
wire n_19039;
wire n_19040;
wire n_19041;
wire n_19042;
wire n_19043;
wire n_19044;
wire n_19045;
wire n_19046;
wire n_19047;
wire n_19048;
wire n_19049;
wire n_19050;
wire n_19051;
wire n_19052;
wire n_19053;
wire n_19054;
wire n_19055;
wire n_19056;
wire n_19057;
wire n_19058;
wire n_19059;
wire n_19060;
wire n_19061;
wire n_19062;
wire n_19063;
wire n_19064;
wire n_19065;
wire n_19066;
wire n_19067;
wire n_19068;
wire n_19069;
wire n_19070;
wire n_19071;
wire n_19072;
wire n_19073;
wire n_19074;
wire n_19075;
wire n_19076;
wire n_19077;
wire n_19078;
wire n_19079;
wire n_19080;
wire n_19081;
wire n_19082;
wire n_19083;
wire n_19084;
wire n_19085;
wire n_19086;
wire n_19087;
wire n_19088;
wire n_19089;
wire n_19090;
wire n_19091;
wire n_19092;
wire n_19093;
wire n_19094;
wire n_19095;
wire n_19096;
wire n_19097;
wire n_19098;
wire n_19099;
wire n_19100;
wire n_19101;
wire n_19102;
wire n_19103;
wire n_19104;
wire n_19105;
wire n_19106;
wire n_19107;
wire n_19108;
wire n_19109;
wire n_19110;
wire n_19111;
wire n_19112;
wire n_19113;
wire n_19114;
wire n_19115;
wire n_19116;
wire n_19117;
wire n_19118;
wire n_19119;
wire n_19120;
wire n_19121;
wire n_19122;
wire n_19123;
wire n_19124;
wire n_19125;
wire n_19126;
wire n_19127;
wire n_19128;
wire n_19129;
wire n_19130;
wire n_19131;
wire n_19132;
wire n_19133;
wire n_19134;
wire n_19135;
wire n_19136;
wire n_19137;
wire n_19138;
wire n_19139;
wire n_19140;
wire n_19141;
wire n_19142;
wire n_19143;
wire n_19144;
wire n_19145;
wire n_19146;
wire n_19147;
wire n_19148;
wire n_19149;
wire n_19150;
wire n_19151;
wire n_19152;
wire n_19153;
wire n_19154;
wire n_19155;
wire n_19156;
wire n_19157;
wire n_19158;
wire n_19159;
wire n_19160;
wire n_19161;
wire n_19162;
wire n_19163;
wire n_19164;
wire n_19165;
wire n_19166;
wire n_19167;
wire n_19168;
wire n_19169;
wire n_19170;
wire n_19171;
wire n_19172;
wire n_19173;
wire n_19174;
wire n_19175;
wire n_19176;
wire n_19177;
wire n_19178;
wire n_19179;
wire n_19180;
wire n_19181;
wire n_19182;
wire n_19183;
wire n_19184;
wire n_19185;
wire n_19186;
wire n_19187;
wire n_19188;
wire n_19189;
wire n_19190;
wire n_19191;
wire n_19192;
wire n_19193;
wire n_19194;
wire n_19195;
wire n_19196;
wire n_19197;
wire n_19198;
wire n_19199;
wire n_19200;
wire n_19201;
wire n_19202;
wire n_19203;
wire n_19204;
wire n_19205;
wire n_19206;
wire n_19207;
wire n_19208;
wire n_19209;
wire n_19210;
wire n_19211;
wire n_19212;
wire n_19213;
wire n_19214;
wire n_19215;
wire n_19216;
wire n_19217;
wire n_19218;
wire n_19219;
wire n_19220;
wire n_19221;
wire n_19222;
wire n_19223;
wire n_19224;
wire n_19225;
wire n_19226;
wire n_19227;
wire n_19228;
wire n_19229;
wire n_19230;
wire n_19231;
wire n_19232;
wire n_19233;
wire n_19234;
wire n_19235;
wire n_19236;
wire n_19237;
wire n_19238;
wire n_19239;
wire n_19240;
wire n_19241;
wire n_19242;
wire n_19243;
wire n_19244;
wire n_19245;
wire n_19246;
wire n_19247;
wire n_19248;
wire n_19249;
wire n_19250;
wire n_19251;
wire n_19252;
wire n_19253;
wire n_19254;
wire n_19255;
wire n_19256;
wire n_19257;
wire n_19258;
wire n_19259;
wire n_19260;
wire n_19261;
wire n_19262;
wire n_19263;
wire n_19264;
wire n_19265;
wire n_19266;
wire n_19267;
wire n_19268;
wire n_19269;
wire n_19270;
wire n_19271;
wire n_19272;
wire n_19273;
wire n_19274;
wire n_19275;
wire n_19276;
wire n_19277;
wire n_19278;
wire n_19279;
wire n_19280;
wire n_19281;
wire n_19282;
wire n_19283;
wire n_19284;
wire n_19285;
wire n_19286;
wire n_19287;
wire n_19288;
wire n_19289;
wire n_19290;
wire n_19291;
wire n_19292;
wire n_19293;
wire n_19294;
wire n_19295;
wire n_19296;
wire n_19297;
wire n_19298;
wire n_19299;
wire n_19300;
wire n_19301;
wire n_19302;
wire n_19303;
wire n_19304;
wire n_19305;
wire n_19306;
wire n_19307;
wire n_19308;
wire n_19309;
wire n_19310;
wire n_19311;
wire n_19312;
wire n_19313;
wire n_19314;
wire n_19315;
wire n_19316;
wire n_19317;
wire n_19318;
wire n_19319;
wire n_19320;
wire n_19321;
wire n_19322;
wire n_19323;
wire n_19324;
wire n_19325;
wire n_19326;
wire n_19327;
wire n_19328;
wire n_19329;
wire n_19330;
wire n_19331;
wire n_19332;
wire n_19333;
wire n_19334;
wire n_19335;
wire n_19336;
wire n_19337;
wire n_19338;
wire n_19339;
wire n_19340;
wire n_19341;
wire n_19342;
wire n_19343;
wire n_19344;
wire n_19345;
wire n_19346;
wire n_19347;
wire n_19348;
wire n_19349;
wire n_19350;
wire n_19351;
wire n_19352;
wire n_19353;
wire n_19354;
wire n_19355;
wire n_19356;
wire n_19357;
wire n_19358;
wire n_19359;
wire n_19360;
wire n_19361;
wire n_19362;
wire n_19363;
wire n_19364;
wire n_19365;
wire n_19366;
wire n_19367;
wire n_19368;
wire n_19369;
wire n_19370;
wire n_19371;
wire n_19372;
wire n_19373;
wire n_19374;
wire n_19375;
wire n_19376;
wire n_19377;
wire n_19378;
wire n_19379;
wire n_19380;
wire n_19381;
wire n_19382;
wire n_19383;
wire n_19384;
wire n_19385;
wire n_19386;
wire n_19387;
wire n_19388;
wire n_19389;
wire n_19390;
wire n_19391;
wire n_19392;
wire n_19393;
wire n_19394;
wire n_19395;
wire n_19396;
wire n_19397;
wire n_19398;
wire n_19399;
wire n_19400;
wire n_19401;
wire n_19402;
wire n_19403;
wire n_19404;
wire n_19405;
wire n_19406;
wire n_19407;
wire n_19408;
wire n_19409;
wire n_19410;
wire n_19411;
wire n_19412;
wire n_19413;
wire n_19414;
wire n_19415;
wire n_19416;
wire n_19417;
wire n_19418;
wire n_19419;
wire n_19420;
wire n_19421;
wire n_19422;
wire n_19423;
wire n_19424;
wire n_19425;
wire n_19426;
wire n_19427;
wire n_19428;
wire n_19429;
wire n_19430;
wire n_19431;
wire n_19432;
wire n_19433;
wire n_19434;
wire n_19435;
wire n_19436;
wire n_19437;
wire n_19438;
wire n_19439;
wire n_19440;
wire n_19441;
wire n_19442;
wire n_19443;
wire n_19444;
wire n_19445;
wire n_19446;
wire n_19447;
wire n_19448;
wire n_19449;
wire n_19450;
wire n_19451;
wire n_19452;
wire n_19453;
wire n_19454;
wire n_19455;
wire n_19456;
wire n_19457;
wire n_19458;
wire n_19459;
wire n_19460;
wire n_19461;
wire n_19462;
wire n_19463;
wire n_19464;
wire n_19465;
wire n_19466;
wire n_19467;
wire n_19468;
wire n_19469;
wire n_19470;
wire n_19471;
wire n_19472;
wire n_19473;
wire n_19474;
wire n_19475;
wire n_19476;
wire n_19477;
wire n_19478;
wire n_19479;
wire n_19480;
wire n_19481;
wire n_19482;
wire n_19483;
wire n_19484;
wire n_19485;
wire n_19486;
wire n_19487;
wire n_19488;
wire n_19489;
wire n_19490;
wire n_19491;
wire n_19492;
wire n_19493;
wire n_19494;
wire n_19495;
wire n_19496;
wire n_19497;
wire n_19498;
wire n_19499;
wire n_19500;
wire n_19501;
wire n_19502;
wire n_19503;
wire n_19504;
wire n_19505;
wire n_19506;
wire n_19507;
wire n_19508;
wire n_19509;
wire n_19510;
wire n_19511;
wire n_19512;
wire n_19513;
wire n_19514;
wire n_19515;
wire n_19516;
wire n_19517;
wire n_19518;
wire n_19519;
wire n_19520;
wire n_19521;
wire n_19522;
wire n_19523;
wire n_19524;
wire n_19525;
wire n_19526;
wire n_19527;
wire n_19528;
wire n_19529;
wire n_19530;
wire n_19531;
wire n_19532;
wire n_19533;
wire n_19534;
wire n_19535;
wire n_19536;
wire n_19537;
wire n_19538;
wire n_19539;
wire n_19540;
wire n_19541;
wire n_19542;
wire n_19543;
wire n_19544;
wire n_19545;
wire n_19546;
wire n_19547;
wire n_19548;
wire n_19549;
wire n_19550;
wire n_19551;
wire n_19552;
wire n_19553;
wire n_19554;
wire n_19555;
wire n_19556;
wire n_19557;
wire n_19558;
wire n_19559;
wire n_19560;
wire n_19561;
wire n_19562;
wire n_19563;
wire n_19564;
wire n_19565;
wire n_19566;
wire n_19567;
wire n_19568;
wire n_19569;
wire n_19570;
wire n_19571;
wire n_19572;
wire n_19573;
wire n_19574;
wire n_19575;
wire n_19576;
wire n_19577;
wire n_19578;
wire n_19579;
wire n_19580;
wire n_19581;
wire n_19582;
wire n_19583;
wire n_19584;
wire n_19585;
wire n_19586;
wire n_19587;
wire n_19588;
wire n_19589;
wire n_19590;
wire n_19591;
wire n_19592;
wire n_19593;
wire n_19594;
wire n_19595;
wire n_19596;
wire n_19597;
wire n_19598;
wire n_19599;
wire n_19600;
wire n_19601;
wire n_19602;
wire n_19603;
wire n_19604;
wire n_19605;
wire n_19606;
wire n_19607;
wire n_19608;
wire n_19609;
wire n_19610;
wire n_19611;
wire n_19612;
wire n_19613;
wire n_19614;
wire n_19615;
wire n_19616;
wire n_19617;
wire n_19618;
wire n_19619;
wire n_19620;
wire n_19621;
wire n_19622;
wire n_19623;
wire n_19624;
wire n_19625;
wire n_19626;
wire n_19627;
wire n_19628;
wire n_19629;
wire n_19630;
wire n_19631;
wire n_19632;
wire n_19633;
wire n_19634;
wire n_19635;
wire n_19636;
wire n_19637;
wire n_19638;
wire n_19639;
wire n_19640;
wire n_19641;
wire n_19642;
wire n_19643;
wire n_19644;
wire n_19645;
wire n_19646;
wire n_19647;
wire n_19648;
wire n_19649;
wire n_19650;
wire n_19651;
wire n_19652;
wire n_19653;
wire n_19654;
wire n_19655;
wire n_19656;
wire n_19657;
wire n_19658;
wire n_19659;
wire n_19660;
wire n_19661;
wire n_19662;
wire n_19663;
wire n_19664;
wire n_19665;
wire n_19666;
wire n_19667;
wire n_19668;
wire n_19669;
wire n_19670;
wire n_19671;
wire n_19672;
wire n_19673;
wire n_19674;
wire n_19675;
wire n_19676;
wire n_19677;
wire n_19678;
wire n_19679;
wire n_19680;
wire n_19681;
wire n_19682;
wire n_19683;
wire n_19684;
wire n_19685;
wire n_19686;
wire n_19687;
wire n_19688;
wire n_19689;
wire n_19690;
wire n_19691;
wire n_19692;
wire n_19693;
wire n_19694;
wire n_19695;
wire n_19696;
wire n_19697;
wire n_19698;
wire n_19699;
wire n_19700;
wire n_19701;
wire n_19702;
wire n_19703;
wire n_19704;
wire n_19705;
wire n_19706;
wire n_19707;
wire n_19708;
wire n_19709;
wire n_19710;
wire n_19711;
wire n_19712;
wire n_19713;
wire n_19714;
wire n_19715;
wire n_19716;
wire n_19717;
wire n_19718;
wire n_19719;
wire n_19720;
wire n_19721;
wire n_19722;
wire n_19723;
wire n_19724;
wire n_19725;
wire n_19726;
wire n_19727;
wire n_19728;
wire n_19729;
wire n_19730;
wire n_19731;
wire n_19732;
wire n_19733;
wire n_19734;
wire n_19735;
wire n_19736;
wire n_19737;
wire n_19738;
wire n_19739;
wire n_19740;
wire n_19741;
wire n_19742;
wire n_19743;
wire n_19744;
wire n_19745;
wire n_19746;
wire n_19747;
wire n_19748;
wire n_19749;
wire n_19750;
wire n_19751;
wire n_19752;
wire n_19753;
wire n_19754;
wire n_19755;
wire n_19756;
wire n_19757;
wire n_19758;
wire n_19759;
wire n_19760;
wire n_19761;
wire n_19762;
wire n_19763;
wire n_19764;
wire n_19765;
wire n_19766;
wire n_19767;
wire n_19768;
wire n_19769;
wire n_19770;
wire n_19771;
wire n_19772;
wire n_19773;
wire n_19774;
wire n_19775;
wire n_19776;
wire n_19777;
wire n_19778;
wire n_19779;
wire n_19780;
wire n_19781;
wire n_19782;
wire n_19783;
wire n_19784;
wire n_19785;
wire n_19786;
wire n_19787;
wire n_19788;
wire n_19789;
wire n_19790;
wire n_19791;
wire n_19792;
wire n_19793;
wire n_19794;
wire n_19795;
wire n_19796;
wire n_19797;
wire n_19798;
wire n_19799;
wire n_19800;
wire n_19801;
wire n_19802;
wire n_19803;
wire n_19804;
wire n_19805;
wire n_19806;
wire n_19807;
wire n_19808;
wire n_19809;
wire n_19810;
wire n_19811;
wire n_19812;
wire n_19813;
wire n_19814;
wire n_19815;
wire n_19816;
wire n_19817;
wire n_19818;
wire n_19819;
wire n_19820;
wire n_19821;
wire n_19822;
wire n_19823;
wire n_19824;
wire n_19825;
wire n_19826;
wire n_19827;
wire n_19828;
wire n_19829;
wire n_19830;
wire n_19831;
wire n_19832;
wire n_19833;
wire n_19834;
wire n_19835;
wire n_19836;
wire n_19837;
wire n_19838;
wire n_19839;
wire n_19840;
wire n_19841;
wire n_19842;
wire n_19843;
wire n_19844;
wire n_19845;
wire n_19846;
wire n_19847;
wire n_19848;
wire n_19849;
wire n_19850;
wire n_19851;
wire n_19852;
wire n_19853;
wire n_19854;
wire n_19855;
wire n_19856;
wire n_19857;
wire n_19858;
wire n_19859;
wire n_19860;
wire n_19861;
wire n_19862;
wire n_19863;
wire n_19864;
wire n_19865;
wire n_19866;
wire n_19867;
wire n_19868;
wire n_19869;
wire n_19870;
wire n_19871;
wire n_19872;
wire n_19873;
wire n_19874;
wire n_19875;
wire n_19876;
wire n_19877;
wire n_19878;
wire n_19879;
wire n_19880;
wire n_19881;
wire n_19882;
wire n_19883;
wire n_19884;
wire n_19885;
wire n_19886;
wire n_19887;
wire n_19888;
wire n_19889;
wire n_19890;
wire n_19891;
wire n_19892;
wire n_19893;
wire n_19894;
wire n_19895;
wire n_19896;
wire n_19897;
wire n_19898;
wire n_19899;
wire n_19900;
wire n_19901;
wire n_19902;
wire n_19903;
wire n_19904;
wire n_19905;
wire n_19906;
wire n_19907;
wire n_19908;
wire n_19909;
wire n_19910;
wire n_19911;
wire n_19912;
wire n_19913;
wire n_19914;
wire n_19915;
wire n_19916;
wire n_19917;
wire n_19918;
wire n_19919;
wire n_19920;
wire n_19921;
wire n_19922;
wire n_19923;
wire n_19924;
wire n_19925;
wire n_19926;
wire n_19927;
wire n_19928;
wire n_19929;
wire n_19930;
wire n_19931;
wire n_19932;
wire n_19933;
wire n_19934;
wire n_19935;
wire n_19936;
wire n_19937;
wire n_19938;
wire n_19939;
wire n_19940;
wire n_19941;
wire n_19942;
wire n_19943;
wire n_19944;
wire n_19945;
wire n_19946;
wire n_19947;
wire n_19948;
wire n_19949;
wire n_19950;
wire n_19951;
wire n_19952;
wire n_19953;
wire n_19954;
wire n_19955;
wire n_19956;
wire n_19957;
wire n_19958;
wire n_19959;
wire n_19960;
wire n_19961;
wire n_19962;
wire n_19963;
wire n_19964;
wire n_19965;
wire n_19966;
wire n_19967;
wire n_19968;
wire n_19969;
wire n_19970;
wire n_19971;
wire n_19972;
wire n_19973;
wire n_19974;
wire n_19975;
wire n_19976;
wire n_19977;
wire n_19978;
wire n_19979;
wire n_19980;
wire n_19981;
wire n_19982;
wire n_19983;
wire n_19984;
wire n_19985;
wire n_19986;
wire n_19987;
wire n_19988;
wire n_19989;
wire n_19990;
wire n_19991;
wire n_19992;
wire n_19993;
wire n_19994;
wire n_19995;
wire n_19996;
wire n_19997;
wire n_19998;
wire n_19999;
wire n_20000;
wire n_20001;
wire n_20002;
wire n_20003;
wire n_20004;
wire n_20005;
wire n_20006;
wire n_20007;
wire n_20008;
wire n_20009;
wire n_20010;
wire n_20011;
wire n_20012;
wire n_20013;
wire n_20014;
wire n_20015;
wire n_20016;
wire n_20017;
wire n_20018;
wire n_20019;
wire n_20020;
wire n_20021;
wire n_20022;
wire n_20023;
wire n_20024;
wire n_20025;
wire n_20026;
wire n_20027;
wire n_20028;
wire n_20029;
wire n_20030;
wire n_20031;
wire n_20032;
wire n_20033;
wire n_20034;
wire n_20035;
wire n_20036;
wire n_20037;
wire n_20038;
wire n_20039;
wire n_20040;
wire n_20041;
wire n_20042;
wire n_20043;
wire n_20044;
wire n_20045;
wire n_20046;
wire n_20047;
wire n_20048;
wire n_20049;
wire n_20050;
wire n_20051;
wire n_20052;
wire n_20053;
wire n_20054;
wire n_20055;
wire n_20056;
wire n_20057;
wire n_20058;
wire n_20059;
wire n_20060;
wire n_20061;
wire n_20062;
wire n_20063;
wire n_20064;
wire n_20065;
wire n_20066;
wire n_20067;
wire n_20068;
wire n_20069;
wire n_20070;
wire n_20071;
wire n_20072;
wire n_20073;
wire n_20074;
wire n_20075;
wire n_20076;
wire n_20077;
wire n_20078;
wire n_20079;
wire n_20080;
wire n_20081;
wire n_20082;
wire n_20083;
wire n_20084;
wire n_20085;
wire n_20086;
wire n_20087;
wire n_20088;
wire n_20089;
wire n_20090;
wire n_20091;
wire n_20092;
wire n_20093;
wire n_20094;
wire n_20095;
wire n_20096;
wire n_20097;
wire n_20098;
wire n_20099;
wire n_20100;
wire n_20101;
wire n_20102;
wire n_20103;
wire n_20104;
wire n_20105;
wire n_20106;
wire n_20107;
wire n_20108;
wire n_20109;
wire n_20110;
wire n_20111;
wire n_20112;
wire n_20113;
wire n_20114;
wire n_20115;
wire n_20116;
wire n_20117;
wire n_20118;
wire n_20119;
wire n_20120;
wire n_20121;
wire n_20122;
wire n_20123;
wire n_20124;
wire n_20125;
wire n_20126;
wire n_20127;
wire n_20128;
wire n_20129;
wire n_20130;
wire n_20131;
wire n_20132;
wire n_20133;
wire n_20134;
wire n_20135;
wire n_20136;
wire n_20137;
wire n_20138;
wire n_20139;
wire n_20140;
wire n_20141;
wire n_20142;
wire n_20143;
wire n_20144;
wire n_20145;
wire n_20146;
wire n_20147;
wire n_20148;
wire n_20149;
wire n_20150;
wire n_20151;
wire n_20152;
wire n_20153;
wire n_20154;
wire n_20155;
wire n_20156;
wire n_20157;
wire n_20158;
wire n_20159;
wire n_20160;
wire n_20161;
wire n_20162;
wire n_20163;
wire n_20164;
wire n_20165;
wire n_20166;
wire n_20167;
wire n_20168;
wire n_20169;
wire n_20170;
wire n_20171;
wire n_20172;
wire n_20173;
wire n_20174;
wire n_20175;
wire n_20176;
wire n_20177;
wire n_20178;
wire n_20179;
wire n_20180;
wire n_20181;
wire n_20182;
wire n_20183;
wire n_20184;
wire n_20185;
wire n_20186;
wire n_20187;
wire n_20188;
wire n_20189;
wire n_20190;
wire n_20191;
wire n_20192;
wire n_20193;
wire n_20194;
wire n_20195;
wire n_20196;
wire n_20197;
wire n_20198;
wire n_20199;
wire n_20200;
wire n_20201;
wire n_20202;
wire n_20203;
wire n_20204;
wire n_20205;
wire n_20206;
wire n_20207;
wire n_20208;
wire n_20209;
wire n_20210;
wire n_20211;
wire n_20212;
wire n_20213;
wire n_20214;
wire n_20215;
wire n_20216;
wire n_20217;
wire n_20218;
wire n_20219;
wire n_20220;
wire n_20221;
wire n_20222;
wire n_20223;
wire n_20224;
wire n_20225;
wire n_20226;
wire n_20227;
wire n_20228;
wire n_20229;
wire n_20230;
wire n_20231;
wire n_20232;
wire n_20233;
wire n_20234;
wire n_20235;
wire n_20236;
wire n_20237;
wire n_20238;
wire n_20239;
wire n_20240;
wire n_20241;
wire n_20242;
wire n_20243;
wire n_20244;
wire n_20245;
wire n_20246;
wire n_20247;
wire n_20248;
wire n_20249;
wire n_20250;
wire n_20251;
wire n_20252;
wire n_20253;
wire n_20254;
wire n_20255;
wire n_20256;
wire n_20257;
wire n_20258;
wire n_20259;
wire n_20260;
wire n_20261;
wire n_20262;
wire n_20263;
wire n_20264;
wire n_20265;
wire n_20266;
wire n_20267;
wire n_20268;
wire n_20269;
wire n_20270;
wire n_20271;
wire n_20272;
wire n_20273;
wire n_20274;
wire n_20275;
wire n_20276;
wire n_20277;
wire n_20278;
wire n_20279;
wire n_20280;
wire n_20281;
wire n_20282;
wire n_20283;
wire n_20284;
wire n_20285;
wire n_20286;
wire n_20287;
wire n_20288;
wire n_20289;
wire n_20290;
wire n_20291;
wire n_20292;
wire n_20293;
wire n_20294;
wire n_20295;
wire n_20296;
wire n_20297;
wire n_20298;
wire n_20299;
wire n_20300;
wire n_20301;
wire n_20302;
wire n_20303;
wire n_20304;
wire n_20305;
wire n_20306;
wire n_20307;
wire n_20308;
wire n_20309;
wire n_20310;
wire n_20311;
wire n_20312;
wire n_20313;
wire n_20314;
wire n_20315;
wire n_20316;
wire n_20317;
wire n_20318;
wire n_20319;
wire n_20320;
wire n_20321;
wire n_20322;
wire n_20323;
wire n_20324;
wire n_20325;
wire n_20326;
wire n_20327;
wire n_20328;
wire n_20329;
wire n_20330;
wire n_20331;
wire n_20332;
wire n_20333;
wire n_20334;
wire n_20335;
wire n_20336;
wire n_20337;
wire n_20338;
wire n_20339;
wire n_20340;
wire n_20341;
wire n_20342;
wire n_20343;
wire n_20344;
wire n_20345;
wire n_20346;
wire n_20347;
wire n_20348;
wire n_20349;
wire n_20350;
wire n_20351;
wire n_20352;
wire n_20353;
wire n_20354;
wire n_20355;
wire n_20356;
wire n_20357;
wire n_20358;
wire n_20359;
wire n_20360;
wire n_20361;
wire n_20362;
wire n_20363;
wire n_20364;
wire n_20365;
wire n_20366;
wire n_20367;
wire n_20368;
wire n_20369;
wire n_20370;
wire n_20371;
wire n_20372;
wire n_20373;
wire n_20374;
wire n_20375;
wire n_20376;
wire n_20377;
wire n_20378;
wire n_20379;
wire n_20380;
wire n_20381;
wire n_20382;
wire n_20383;
wire n_20384;
wire n_20385;
wire n_20386;
wire n_20387;
wire n_20388;
wire n_20389;
wire n_20390;
wire n_20391;
wire n_20392;
wire n_20393;
wire n_20394;
wire n_20395;
wire n_20396;
wire n_20397;
wire n_20398;
wire n_20399;
wire n_20400;
wire n_20401;
wire n_20402;
wire n_20403;
wire n_20404;
wire n_20405;
wire n_20406;
wire n_20407;
wire n_20408;
wire n_20409;
wire n_20410;
wire n_20411;
wire n_20412;
wire n_20413;
wire n_20414;
wire n_20415;
wire n_20416;
wire n_20417;
wire n_20418;
wire n_20419;
wire n_20420;
wire n_20421;
wire n_20422;
wire n_20423;
wire n_20424;
wire n_20425;
wire n_20426;
wire n_20427;
wire n_20428;
wire n_20429;
wire n_20430;
wire n_20431;
wire n_20432;
wire n_20433;
wire n_20434;
wire n_20435;
wire n_20436;
wire n_20437;
wire n_20438;
wire n_20439;
wire n_20440;
wire n_20441;
wire n_20442;
wire n_20443;
wire n_20444;
wire n_20445;
wire n_20446;
wire n_20447;
wire n_20448;
wire n_20449;
wire n_20450;
wire n_20451;
wire n_20452;
wire n_20453;
wire n_20454;
wire n_20455;
wire n_20456;
wire n_20457;
wire n_20458;
wire n_20459;
wire n_20460;
wire n_20461;
wire n_20462;
wire n_20463;
wire n_20464;
wire n_20465;
wire n_20466;
wire n_20467;
wire n_20468;
wire n_20469;
wire n_20470;
wire n_20471;
wire n_20472;
wire n_20473;
wire n_20474;
wire n_20475;
wire n_20476;
wire n_20477;
wire n_20478;
wire n_20479;
wire n_20480;
wire n_20481;
wire n_20482;
wire n_20483;
wire n_20484;
wire n_20485;
wire n_20486;
wire n_20487;
wire n_20488;
wire n_20489;
wire n_20490;
wire n_20491;
wire n_20492;
wire n_20493;
wire n_20494;
wire n_20495;
wire n_20496;
wire n_20497;
wire n_20498;
wire n_20499;
wire n_20500;
wire n_20501;
wire n_20502;
wire n_20503;
wire n_20504;
wire n_20505;
wire n_20506;
wire n_20507;
wire n_20508;
wire n_20509;
wire n_20510;
wire n_20511;
wire n_20512;
wire n_20513;
wire n_20514;
wire n_20515;
wire n_20516;
wire n_20517;
wire n_20518;
wire n_20519;
wire n_20520;
wire n_20521;
wire n_20522;
wire n_20523;
wire n_20524;
wire n_20525;
wire n_20526;
wire n_20527;
wire n_20528;
wire n_20529;
wire n_20530;
wire n_20531;
wire n_20532;
wire n_20533;
wire n_20534;
wire n_20535;
wire n_20536;
wire n_20537;
wire n_20538;
wire n_20539;
wire n_20540;
wire n_20541;
wire n_20542;
wire n_20543;
wire n_20544;
wire n_20545;
wire n_20546;
wire n_20547;
wire n_20548;
wire n_20549;
wire n_20550;
wire n_20551;
wire n_20552;
wire n_20553;
wire n_20554;
wire n_20555;
wire n_20556;
wire n_20557;
wire n_20558;
wire n_20559;
wire n_20560;
wire n_20561;
wire n_20562;
wire n_20563;
wire n_20564;
wire n_20565;
wire n_20566;
wire n_20567;
wire n_20568;
wire n_20569;
wire n_20570;
wire n_20571;
wire n_20572;
wire n_20573;
wire n_20574;
wire n_20575;
wire n_20576;
wire n_20577;
wire n_20578;
wire n_20579;
wire n_20580;
wire n_20581;
wire n_20582;
wire n_20583;
wire n_20584;
wire n_20585;
wire n_20586;
wire n_20587;
wire n_20588;
wire n_20589;
wire n_20590;
wire n_20591;
wire n_20592;
wire n_20593;
wire n_20594;
wire n_20595;
wire n_20596;
wire n_20597;
wire n_20598;
wire n_20599;
wire n_20600;
wire n_20601;
wire n_20602;
wire n_20603;
wire n_20604;
wire n_20605;
wire n_20606;
wire n_20607;
wire n_20608;
wire n_20609;
wire n_20610;
wire n_20611;
wire n_20612;
wire n_20613;
wire n_20614;
wire n_20615;
wire n_20616;
wire n_20617;
wire n_20618;
wire n_20619;
wire n_20620;
wire n_20621;
wire n_20622;
wire n_20623;
wire n_20624;
wire n_20625;
wire n_20626;
wire n_20627;
wire n_20628;
wire n_20629;
wire n_20630;
wire n_20631;
wire n_20632;
wire n_20633;
wire n_20634;
wire n_20635;
wire n_20636;
wire n_20637;
wire n_20638;
wire n_20639;
wire n_20640;
wire n_20641;
wire n_20642;
wire n_20643;
wire n_20644;
wire n_20645;
wire n_20646;
wire n_20647;
wire n_20648;
wire n_20649;
wire n_20650;
wire n_20651;
wire n_20652;
wire n_20653;
wire n_20654;
wire n_20655;
wire n_20656;
wire n_20657;
wire n_20658;
wire n_20659;
wire n_20660;
wire n_20661;
wire n_20662;
wire n_20663;
wire n_20664;
wire n_20665;
wire n_20666;
wire n_20667;
wire n_20668;
wire n_20669;
wire n_20670;
wire n_20671;
wire n_20672;
wire n_20673;
wire n_20674;
wire n_20675;
wire n_20676;
wire n_20677;
wire n_20678;
wire n_20679;
wire n_20680;
wire n_20681;
wire n_20682;
wire n_20683;
wire n_20684;
wire n_20685;
wire n_20686;
wire n_20687;
wire n_20688;
wire n_20689;
wire n_20690;
wire n_20691;
wire n_20692;
wire n_20693;
wire n_20694;
wire n_20695;
wire n_20696;
wire n_20697;
wire n_20698;
wire n_20699;
wire n_20700;
wire n_20701;
wire n_20702;
wire n_20703;
wire n_20704;
wire n_20705;
wire n_20706;
wire n_20707;
wire n_20708;
wire n_20709;
wire n_20710;
wire n_20711;
wire n_20712;
wire n_20713;
wire n_20714;
wire n_20715;
wire n_20716;
wire n_20717;
wire n_20718;
wire n_20719;
wire n_20720;
wire n_20721;
wire n_20722;
wire n_20723;
wire n_20724;
wire n_20725;
wire n_20726;
wire n_20727;
wire n_20728;
wire n_20729;
wire n_20730;
wire n_20731;
wire n_20732;
wire n_20733;
wire n_20734;
wire n_20735;
wire n_20736;
wire n_20737;
wire n_20738;
wire n_20739;
wire n_20740;
wire n_20741;
wire n_20742;
wire n_20743;
wire n_20744;
wire n_20745;
wire n_20746;
wire n_20747;
wire n_20748;
wire n_20749;
wire n_20750;
wire n_20751;
wire n_20752;
wire n_20753;
wire n_20754;
wire n_20755;
wire n_20756;
wire n_20757;
wire n_20758;
wire n_20759;
wire n_20760;
wire n_20761;
wire n_20762;
wire n_20763;
wire n_20764;
wire n_20765;
wire n_20766;
wire n_20767;
wire n_20768;
wire n_20769;
wire n_20770;
wire n_20771;
wire n_20772;
wire n_20773;
wire n_20774;
wire n_20775;
wire n_20776;
wire n_20777;
wire n_20778;
wire n_20779;
wire n_20780;
wire n_20781;
wire n_20782;
wire n_20783;
wire n_20784;
wire n_20785;
wire n_20786;
wire n_20787;
wire n_20788;
wire n_20789;
wire n_20790;
wire n_20791;
wire n_20792;
wire n_20793;
wire n_20794;
wire n_20795;
wire n_20796;
wire n_20797;
wire n_20798;
wire n_20799;
wire n_20800;
wire n_20801;
wire n_20802;
wire n_20803;
wire n_20804;
wire n_20805;
wire n_20806;
wire n_20807;
wire n_20808;
wire n_20809;
wire n_20810;
wire n_20811;
wire n_20812;
wire n_20813;
wire n_20814;
wire n_20815;
wire n_20816;
wire n_20817;
wire n_20818;
wire n_20819;
wire n_20820;
wire n_20821;
wire n_20822;
wire n_20823;
wire n_20824;
wire n_20825;
wire n_20826;
wire n_20827;
wire n_20828;
wire n_20829;
wire n_20830;
wire n_20831;
wire n_20832;
wire n_20833;
wire n_20834;
wire n_20835;
wire n_20836;
wire n_20837;
wire n_20838;
wire n_20839;
wire n_20840;
wire n_20841;
wire n_20842;
wire n_20843;
wire n_20844;
wire n_20845;
wire n_20846;
wire n_20847;
wire n_20848;
wire n_20849;
wire n_20850;
wire n_20851;
wire n_20852;
wire n_20853;
wire n_20854;
wire n_20855;
wire n_20856;
wire n_20857;
wire n_20858;
wire n_20859;
wire n_20860;
wire n_20861;
wire n_20862;
wire n_20863;
wire n_20864;
wire n_20865;
wire n_20866;
wire n_20867;
wire n_20868;
wire n_20869;
wire n_20870;
wire n_20871;
wire n_20872;
wire n_20873;
wire n_20874;
wire n_20875;
wire n_20876;
wire n_20877;
wire n_20878;
wire n_20879;
wire n_20880;
wire n_20881;
wire n_20882;
wire n_20883;
wire n_20884;
wire n_20885;
wire n_20886;
wire n_20887;
wire n_20888;
wire n_20889;
wire n_20890;
wire n_20891;
wire n_20892;
wire n_20893;
wire n_20894;
wire n_20895;
wire n_20896;
wire n_20897;
wire n_20898;
wire n_20899;
wire n_20900;
wire n_20901;
wire n_20902;
wire n_20903;
wire n_20904;
wire n_20905;
wire n_20906;
wire n_20907;
wire n_20908;
wire n_20909;
wire n_20910;
wire n_20911;
wire n_20912;
wire n_20913;
wire n_20914;
wire n_20915;
wire n_20916;
wire n_20917;
wire n_20918;
wire n_20919;
wire n_20920;
wire n_20921;
wire n_20922;
wire n_20923;
wire n_20924;
wire n_20925;
wire n_20926;
wire n_20927;
wire n_20928;
wire n_20929;
wire n_20930;
wire n_20931;
wire n_20932;
wire n_20933;
wire n_20934;
wire n_20935;
wire n_20936;
wire n_20937;
wire n_20938;
wire n_20939;
wire n_20940;
wire n_20941;
wire n_20942;
wire n_20943;
wire n_20944;
wire n_20945;
wire n_20946;
wire n_20947;
wire n_20948;
wire n_20949;
wire n_20950;
wire n_20951;
wire n_20952;
wire n_20953;
wire n_20954;
wire n_20955;
wire n_20956;
wire n_20957;
wire n_20958;
wire n_20959;
wire n_20960;
wire n_20961;
wire n_20962;
wire n_20963;
wire n_20964;
wire n_20965;
wire n_20966;
wire n_20967;
wire n_20968;
wire n_20969;
wire n_20970;
wire n_20971;
wire n_20972;
wire n_20973;
wire n_20974;
wire n_20975;
wire n_20976;
wire n_20977;
wire n_20978;
wire n_20979;
wire n_20980;
wire n_20981;
wire n_20982;
wire n_20983;
wire n_20984;
wire n_20985;
wire n_20986;
wire n_20987;
wire n_20988;
wire n_20989;
wire n_20990;
wire n_20991;
wire n_20992;
wire n_20993;
wire n_20994;
wire n_20995;
wire n_20996;
wire n_20997;
wire n_20998;
wire n_20999;
wire n_21000;
wire n_21001;
wire n_21002;
wire n_21003;
wire n_21004;
wire n_21005;
wire n_21006;
wire n_21007;
wire n_21008;
wire n_21009;
wire n_21010;
wire n_21011;
wire n_21012;
wire n_21013;
wire n_21014;
wire n_21015;
wire n_21016;
wire n_21017;
wire n_21018;
wire n_21019;
wire n_21020;
wire n_21021;
wire n_21022;
wire n_21023;
wire n_21024;
wire n_21025;
wire n_21026;
wire n_21027;
wire n_21028;
wire n_21029;
wire n_21030;
wire n_21031;
wire n_21032;
wire n_21033;
wire n_21034;
wire n_21035;
wire n_21036;
wire n_21037;
wire n_21038;
wire n_21039;
wire n_21040;
wire n_21041;
wire n_21042;
wire n_21043;
wire n_21044;
wire n_21045;
wire n_21046;
wire n_21047;
wire n_21048;
wire n_21049;
wire n_21050;
wire n_21051;
wire n_21052;
wire n_21053;
wire n_21054;
wire n_21055;
wire n_21056;
wire n_21057;
wire n_21058;
wire n_21059;
wire n_21060;
wire n_21061;
wire n_21062;
wire n_21063;
wire n_21064;
wire n_21065;
wire n_21066;
wire n_21067;
wire n_21068;
wire n_21069;
wire n_21070;
wire n_21071;
wire n_21072;
wire n_21073;
wire n_21074;
wire n_21075;
wire n_21076;
wire n_21077;
wire n_21078;
wire n_21079;
wire n_21080;
wire n_21081;
wire n_21082;
wire n_21083;
wire n_21084;
wire n_21085;
wire n_21086;
wire n_21087;
wire n_21088;
wire n_21089;
wire n_21090;
wire n_21091;
wire n_21092;
wire n_21093;
wire n_21094;
wire n_21095;
wire n_21096;
wire n_21097;
wire n_21098;
wire n_21099;
wire n_21100;
wire n_21101;
wire n_21102;
wire n_21103;
wire n_21104;
wire n_21105;
wire n_21106;
wire n_21107;
wire n_21108;
wire n_21109;
wire n_21110;
wire n_21111;
wire n_21112;
wire n_21113;
wire n_21114;
wire n_21115;
wire n_21116;
wire n_21117;
wire n_21118;
wire n_21119;
wire n_21120;
wire n_21121;
wire n_21122;
wire n_21123;
wire n_21124;
wire n_21125;
wire n_21126;
wire n_21127;
wire n_21128;
wire n_21129;
wire n_21130;
wire n_21131;
wire n_21132;
wire n_21133;
wire n_21134;
wire n_21135;
wire n_21136;
wire n_21137;
wire n_21138;
wire n_21139;
wire n_21140;
wire n_21141;
wire n_21142;
wire n_21143;
wire n_21144;
wire n_21145;
wire n_21146;
wire n_21147;
wire n_21148;
wire n_21149;
wire n_21150;
wire n_21151;
wire n_21152;
wire n_21153;
wire n_21154;
wire n_21155;
wire n_21156;
wire n_21157;
wire n_21158;
wire n_21159;
wire n_21160;
wire n_21161;
wire n_21162;
wire n_21163;
wire n_21164;
wire n_21165;
wire n_21166;
wire n_21167;
wire n_21168;
wire n_21169;
wire n_21170;
wire n_21171;
wire n_21172;
wire n_21173;
wire n_21174;
wire n_21175;
wire n_21176;
wire n_21177;
wire n_21178;
wire n_21179;
wire n_21180;
wire n_21181;
wire n_21182;
wire n_21183;
wire n_21184;
wire n_21185;
wire n_21186;
wire n_21187;
wire n_21188;
wire n_21189;
wire n_21190;
wire n_21191;
wire n_21192;
wire n_21193;
wire n_21194;
wire n_21195;
wire n_21196;
wire n_21197;
wire n_21198;
wire n_21199;
wire n_21200;
wire n_21201;
wire n_21202;
wire n_21203;
wire n_21204;
wire n_21205;
wire n_21206;
wire n_21207;
wire n_21208;
wire n_21209;
wire n_21210;
wire n_21211;
wire n_21212;
wire n_21213;
wire n_21214;
wire n_21215;
wire n_21216;
wire n_21217;
wire n_21218;
wire n_21219;
wire n_21220;
wire n_21221;
wire n_21222;
wire n_21223;
wire n_21224;
wire n_21225;
wire n_21226;
wire n_21227;
wire n_21228;
wire n_21229;
wire n_21230;
wire n_21231;
wire n_21232;
wire n_21233;
wire n_21234;
wire n_21235;
wire n_21236;
wire n_21237;
wire n_21238;
wire n_21239;
wire n_21240;
wire n_21241;
wire n_21242;
wire n_21243;
wire n_21244;
wire n_21245;
wire n_21246;
wire n_21247;
wire n_21248;
wire n_21249;
wire n_21250;
wire n_21251;
wire n_21252;
wire n_21253;
wire n_21254;
wire n_21255;
wire n_21256;
wire n_21257;
wire n_21258;
wire n_21259;
wire n_21260;
wire n_21261;
wire n_21262;
wire n_21263;
wire n_21264;
wire n_21265;
wire n_21266;
wire n_21267;
wire n_21268;
wire n_21269;
wire n_21270;
wire n_21271;
wire n_21272;
wire n_21273;
wire n_21274;
wire n_21275;
wire n_21276;
wire n_21277;
wire n_21278;
wire n_21279;
wire n_21280;
wire n_21281;
wire n_21282;
wire n_21283;
wire n_21284;
wire n_21285;
wire n_21286;
wire n_21287;
wire n_21288;
wire n_21289;
wire n_21290;
wire n_21291;
wire n_21292;
wire n_21293;
wire n_21294;
wire n_21295;
wire n_21296;
wire n_21297;
wire n_21298;
wire n_21299;
wire n_21300;
wire n_21301;
wire n_21302;
wire n_21303;
wire n_21304;
wire n_21305;
wire n_21306;
wire n_21307;
wire n_21308;
wire n_21309;
wire n_21310;
wire n_21311;
wire n_21312;
wire n_21313;
wire n_21314;
wire n_21315;
wire n_21316;
wire n_21317;
wire n_21318;
wire n_21319;
wire n_21320;
wire n_21321;
wire n_21322;
wire n_21323;
wire n_21324;
wire n_21325;
wire n_21326;
wire n_21327;
wire n_21328;
wire n_21329;
wire n_21330;
wire n_21331;
wire n_21332;
wire n_21333;
wire n_21334;
wire n_21335;
wire n_21336;
wire n_21337;
wire n_21338;
wire n_21339;
wire n_21340;
wire n_21341;
wire n_21342;
wire n_21343;
wire n_21344;
wire n_21345;
wire n_21346;
wire n_21347;
wire n_21348;
wire n_21349;
wire n_21350;
wire n_21351;
wire n_21352;
wire n_21353;
wire n_21354;
wire n_21355;
wire n_21356;
wire n_21357;
wire n_21358;
wire n_21359;
wire n_21360;
wire n_21361;
wire n_21362;
wire n_21363;
wire n_21364;
wire n_21365;
wire n_21366;
wire n_21367;
wire n_21368;
wire n_21369;
wire n_21370;
wire n_21371;
wire n_21372;
wire n_21373;
wire n_21374;
wire n_21375;
wire n_21376;
wire n_21377;
wire n_21378;
wire n_21379;
wire n_21380;
wire n_21381;
wire n_21382;
wire n_21383;
wire n_21384;
wire n_21385;
wire n_21386;
wire n_21387;
wire n_21388;
wire n_21389;
wire n_21390;
wire n_21391;
wire n_21392;
wire n_21393;
wire n_21394;
wire n_21395;
wire n_21396;
wire n_21397;
wire n_21398;
wire n_21399;
wire n_21400;
wire n_21401;
wire n_21402;
wire n_21403;
wire n_21404;
wire n_21405;
wire n_21406;
wire n_21407;
wire n_21408;
wire n_21409;
wire n_21410;
wire n_21411;
wire n_21412;
wire n_21413;
wire n_21414;
wire n_21415;
wire n_21416;
wire n_21417;
wire n_21418;
wire n_21419;
wire n_21420;
wire n_21421;
wire n_21422;
wire n_21423;
wire n_21424;
wire n_21425;
wire n_21426;
wire n_21427;
wire n_21428;
wire n_21429;
wire n_21430;
wire n_21431;
wire n_21432;
wire n_21433;
wire n_21434;
wire n_21435;
wire n_21436;
wire n_21437;
wire n_21438;
wire n_21439;
wire n_21440;
wire n_21441;
wire n_21442;
wire n_21443;
wire n_21444;
wire n_21445;
wire n_21446;
wire n_21447;
wire n_21448;
wire n_21449;
wire n_21450;
wire n_21451;
wire n_21452;
wire n_21453;
wire n_21454;
wire n_21455;
wire n_21456;
wire n_21457;
wire n_21458;
wire n_21459;
wire n_21460;
wire n_21461;
wire n_21462;
wire n_21463;
wire n_21464;
wire n_21465;
wire n_21466;
wire n_21467;
wire n_21468;
wire n_21469;
wire n_21470;
wire n_21471;
wire n_21472;
wire n_21473;
wire n_21474;
wire n_21475;
wire n_21476;
wire n_21477;
wire n_21478;
wire n_21479;
wire n_21480;
wire n_21481;
wire n_21482;
wire n_21483;
wire n_21484;
wire n_21485;
wire n_21486;
wire n_21487;
wire n_21488;
wire n_21489;
wire n_21490;
wire n_21491;
wire n_21492;
wire n_21493;
wire n_21494;
wire n_21495;
wire n_21496;
wire n_21497;
wire n_21498;
wire n_21499;
wire n_21500;
wire n_21501;
wire n_21502;
wire n_21503;
wire n_21504;
wire n_21505;
wire n_21506;
wire n_21507;
wire n_21508;
wire n_21509;
wire n_21510;
wire n_21511;
wire n_21512;
wire n_21513;
wire n_21514;
wire n_21515;
wire n_21516;
wire n_21517;
wire n_21518;
wire n_21519;
wire n_21520;
wire n_21521;
wire n_21522;
wire n_21523;
wire n_21524;
wire n_21525;
wire n_21526;
wire n_21527;
wire n_21528;
wire n_21529;
wire n_21530;
wire n_21531;
wire n_21532;
wire n_21533;
wire n_21534;
wire n_21535;
wire n_21536;
wire n_21537;
wire n_21538;
wire n_21539;
wire n_21540;
wire n_21541;
wire n_21542;
wire n_21543;
wire n_21544;
wire n_21545;
wire n_21546;
wire n_21547;
wire n_21548;
wire n_21549;
wire n_21550;
wire n_21551;
wire n_21552;
wire n_21553;
wire n_21554;
wire n_21555;
wire n_21556;
wire n_21557;
wire n_21558;
wire n_21559;
wire n_21560;
wire n_21561;
wire n_21562;
wire n_21563;
wire n_21564;
wire n_21565;
wire n_21566;
wire n_21567;
wire n_21568;
wire n_21569;
wire n_21570;
wire n_21571;
wire n_21572;
wire n_21573;
wire n_21574;
wire n_21575;
wire n_21576;
wire n_21577;
wire n_21578;
wire n_21579;
wire n_21580;
wire n_21581;
wire n_21582;
wire n_21583;
wire n_21584;
wire n_21585;
wire n_21586;
wire n_21587;
wire n_21588;
wire n_21589;
wire n_21590;
wire n_21591;
wire n_21592;
wire n_21593;
wire n_21594;
wire n_21595;
wire n_21596;
wire n_21597;
wire n_21598;
wire n_21599;
wire n_21600;
wire n_21601;
wire n_21602;
wire n_21603;
wire n_21604;
wire n_21605;
wire n_21606;
wire n_21607;
wire n_21608;
wire n_21609;
wire n_21610;
wire n_21611;
wire n_21612;
wire n_21613;
wire n_21614;
wire n_21615;
wire n_21616;
wire n_21617;
wire n_21618;
wire n_21619;
wire n_21620;
wire n_21621;
wire n_21622;
wire n_21623;
wire n_21624;
wire n_21625;
wire n_21626;
wire n_21627;
wire n_21628;
wire n_21629;
wire n_21630;
wire n_21631;
wire n_21632;
wire n_21633;
wire n_21634;
wire n_21635;
wire n_21636;
wire n_21637;
wire n_21638;
wire n_21639;
wire n_21640;
wire n_21641;
wire n_21642;
wire n_21643;
wire n_21644;
wire n_21645;
wire n_21646;
wire n_21647;
wire n_21648;
wire n_21649;
wire n_21650;
wire n_21651;
wire n_21652;
wire n_21653;
wire n_21654;
wire n_21655;
wire n_21656;
wire n_21657;
wire n_21658;
wire n_21659;
wire n_21660;
wire n_21661;
wire n_21662;
wire n_21663;
wire n_21664;
wire n_21665;
wire n_21666;
wire n_21667;
wire n_21668;
wire n_21669;
wire n_21670;
wire n_21671;
wire n_21672;
wire n_21673;
wire n_21674;
wire n_21675;
wire n_21676;
wire n_21677;
wire n_21678;
wire n_21679;
wire n_21680;
wire n_21681;
wire n_21682;
wire n_21683;
wire n_21684;
wire n_21685;
wire n_21686;
wire n_21687;
wire n_21688;
wire n_21689;
wire n_21690;
wire n_21691;
wire n_21692;
wire n_21693;
wire n_21694;
wire n_21695;
wire n_21696;
wire n_21697;
wire n_21698;
wire n_21699;
wire n_21700;
wire n_21701;
wire n_21702;
wire n_21703;
wire n_21704;
wire n_21705;
wire n_21706;
wire n_21707;
wire n_21708;
wire n_21709;
wire n_21710;
wire n_21711;
wire n_21712;
wire n_21713;
wire n_21714;
wire n_21715;
wire n_21716;
wire n_21717;
wire n_21718;
wire n_21719;
wire n_21720;
wire n_21721;
wire n_21722;
wire n_21723;
wire n_21724;
wire n_21725;
wire n_21726;
wire n_21727;
wire n_21728;
wire n_21729;
wire n_21730;
wire n_21731;
wire n_21732;
wire n_21733;
wire n_21734;
wire n_21735;
wire n_21736;
wire n_21737;
wire n_21738;
wire n_21739;
wire n_21740;
wire n_21741;
wire n_21742;
wire n_21743;
wire n_21744;
wire n_21745;
wire n_21746;
wire n_21747;
wire n_21748;
wire n_21749;
wire n_21750;
wire n_21751;
wire n_21752;
wire n_21753;
wire n_21754;
wire n_21755;
wire n_21756;
wire n_21757;
wire n_21758;
wire n_21759;
wire n_21760;
wire n_21761;
wire n_21762;
wire n_21763;
wire n_21764;
wire n_21765;
wire n_21766;
wire n_21767;
wire n_21768;
wire n_21769;
wire n_21770;
wire n_21771;
wire n_21772;
wire n_21773;
wire n_21774;
wire n_21775;
wire n_21776;
wire n_21777;
wire n_21778;
wire n_21779;
wire n_21780;
wire n_21781;
wire n_21782;
wire n_21783;
wire n_21784;
wire n_21785;
wire n_21786;
wire n_21787;
wire n_21788;
wire n_21789;
wire n_21790;
wire n_21791;
wire n_21792;
wire n_21793;
wire n_21794;
wire n_21795;
wire n_21796;
wire n_21797;
wire n_21798;
wire n_21799;
wire n_21800;
wire n_21801;
wire n_21802;
wire n_21803;
wire n_21804;
wire n_21805;
wire n_21806;
wire n_21807;
wire n_21808;
wire n_21809;
wire n_21810;
wire n_21811;
wire n_21812;
wire n_21813;
wire n_21814;
wire n_21815;
wire n_21816;
wire n_21817;
wire n_21818;
wire n_21819;
wire n_21820;
wire n_21821;
wire n_21822;
wire n_21823;
wire n_21824;
wire n_21825;
wire n_21826;
wire n_21827;
wire n_21828;
wire n_21829;
wire n_21830;
wire n_21831;
wire n_21832;
wire n_21833;
wire n_21834;
wire n_21835;
wire n_21836;
wire n_21837;
wire n_21838;
wire n_21839;
wire n_21840;
wire n_21841;
wire n_21842;
wire n_21843;
wire n_21844;
wire n_21845;
wire n_21846;
wire n_21847;
wire n_21848;
wire n_21849;
wire n_21850;
wire n_21851;
wire n_21852;
wire n_21853;
wire n_21854;
wire n_21855;
wire n_21856;
wire n_21857;
wire n_21858;
wire n_21859;
wire n_21860;
wire n_21861;
wire n_21862;
wire n_21863;
wire n_21864;
wire n_21865;
wire n_21866;
wire n_21867;
wire n_21868;
wire n_21869;
wire n_21870;
wire n_21871;
wire n_21872;
wire n_21873;
wire n_21874;
wire n_21875;
wire n_21876;
wire n_21877;
wire n_21878;
wire n_21879;
wire n_21880;
wire n_21881;
wire n_21882;
wire n_21883;
wire n_21884;
wire n_21885;
wire n_21886;
wire n_21887;
wire n_21888;
wire n_21889;
wire n_21890;
wire n_21891;
wire n_21892;
wire n_21893;
wire n_21894;
wire n_21895;
wire n_21896;
wire n_21897;
wire n_21898;
wire n_21899;
wire n_21900;
wire n_21901;
wire n_21902;
wire n_21903;
wire n_21904;
wire n_21905;
wire n_21906;
wire n_21907;
wire n_21908;
wire n_21909;
wire n_21910;
wire n_21911;
wire n_21912;
wire n_21913;
wire n_21914;
wire n_21915;
wire n_21916;
wire n_21917;
wire n_21918;
wire n_21919;
wire n_21920;
wire n_21921;
wire n_21922;
wire n_21923;
wire n_21924;
wire n_21925;
wire n_21926;
wire n_21927;
wire n_21928;
wire n_21929;
wire n_21930;
wire n_21931;
wire n_21932;
wire n_21933;
wire n_21934;
wire n_21935;
wire n_21936;
wire n_21937;
wire n_21938;
wire n_21939;
wire n_21940;
wire n_21941;
wire n_21942;
wire n_21943;
wire n_21944;
wire n_21945;
wire n_21946;
wire n_21947;
wire n_21948;
wire n_21949;
wire n_21950;
wire n_21951;
wire n_21952;
wire n_21953;
wire n_21954;
wire n_21955;
wire n_21956;
wire n_21957;
wire n_21958;
wire n_21959;
wire n_21960;
wire n_21961;
wire n_21962;
wire n_21963;
wire n_21964;
wire n_21965;
wire n_21966;
wire n_21967;
wire n_21968;
wire n_21969;
wire n_21970;
wire n_21971;
wire n_21972;
wire n_21973;
wire n_21974;
wire n_21975;
wire n_21976;
wire n_21977;
wire n_21978;
wire n_21979;
wire n_21980;
wire n_21981;
wire n_21982;
wire n_21983;
wire n_21984;
wire n_21985;
wire n_21986;
wire n_21987;
wire n_21988;
wire n_21989;
wire n_21990;
wire n_21991;
wire n_21992;
wire n_21993;
wire n_21994;
wire n_21995;
wire n_21996;
wire n_21997;
wire n_21998;
wire n_21999;
wire n_22000;
wire n_22001;
wire n_22002;
wire n_22003;
wire n_22004;
wire n_22005;
wire n_22006;
wire n_22007;
wire n_22008;
wire n_22009;
wire n_22010;
wire n_22011;
wire n_22012;
wire n_22013;
wire n_22014;
wire n_22015;
wire n_22016;
wire n_22017;
wire n_22018;
wire n_22019;
wire n_22020;
wire n_22021;
wire n_22022;
wire n_22023;
wire n_22024;
wire n_22025;
wire n_22026;
wire n_22027;
wire n_22028;
wire n_22029;
wire n_22030;
wire n_22031;
wire n_22032;
wire n_22033;
wire n_22034;
wire n_22035;
wire n_22036;
wire n_22037;
wire n_22038;
wire n_22039;
wire n_22040;
wire n_22041;
wire n_22042;
wire n_22043;
wire n_22044;
wire n_22045;
wire n_22046;
wire n_22047;
wire n_22048;
wire n_22049;
wire n_22050;
wire n_22051;
wire n_22052;
wire n_22053;
wire n_22054;
wire n_22055;
wire n_22056;
wire n_22057;
wire n_22058;
wire n_22059;
wire n_22060;
wire n_22061;
wire n_22062;
wire n_22063;
wire n_22064;
wire n_22065;
wire n_22066;
wire n_22067;
wire n_22068;
wire n_22069;
wire n_22070;
wire n_22071;
wire n_22072;
wire n_22073;
wire n_22074;
wire n_22075;
wire n_22076;
wire n_22077;
wire n_22078;
wire n_22079;
wire n_22080;
wire n_22081;
wire n_22082;
wire n_22083;
wire n_22084;
wire n_22085;
wire n_22086;
wire n_22087;
wire n_22088;
wire n_22089;
wire n_22090;
wire n_22091;
wire n_22092;
wire n_22093;
wire n_22094;
wire n_22095;
wire n_22096;
wire n_22097;
wire n_22098;
wire n_22099;
wire n_22100;
wire n_22101;
wire n_22102;
wire n_22103;
wire n_22104;
wire n_22105;
wire n_22106;
wire n_22107;
wire n_22108;
wire n_22109;
wire n_22110;
wire n_22111;
wire n_22112;
wire n_22113;
wire n_22114;
wire n_22115;
wire n_22116;
wire n_22117;
wire n_22118;
wire n_22119;
wire n_22120;
wire n_22121;
wire n_22122;
wire n_22123;
wire n_22124;
wire n_22125;
wire n_22126;
wire n_22127;
wire n_22128;
wire n_22129;
wire n_22130;
wire n_22131;
wire n_22132;
wire n_22133;
wire n_22134;
wire n_22135;
wire n_22136;
wire n_22137;
wire n_22138;
wire n_22139;
wire n_22140;
wire n_22141;
wire n_22142;
wire n_22143;
wire n_22144;
wire n_22145;
wire n_22146;
wire n_22147;
wire n_22148;
wire n_22149;
wire n_22150;
wire n_22151;
wire n_22152;
wire n_22153;
wire n_22154;
wire n_22155;
wire n_22156;
wire n_22157;
wire n_22158;
wire n_22159;
wire n_22160;
wire n_22161;
wire n_22162;
wire n_22163;
wire n_22164;
wire n_22165;
wire n_22166;
wire n_22167;
wire n_22168;
wire n_22169;
wire n_22170;
wire n_22171;
wire n_22172;
wire n_22173;
wire n_22174;
wire n_22175;
wire n_22176;
wire n_22177;
wire n_22178;
wire n_22179;
wire n_22180;
wire n_22181;
wire n_22182;
wire n_22183;
wire n_22184;
wire n_22185;
wire n_22186;
wire n_22187;
wire n_22188;
wire n_22189;
wire n_22190;
wire n_22191;
wire n_22192;
wire n_22193;
wire n_22194;
wire n_22195;
wire n_22196;
wire n_22197;
wire n_22198;
wire n_22199;
wire n_22200;
wire n_22201;
wire n_22202;
wire n_22203;
wire n_22204;
wire n_22205;
wire n_22206;
wire n_22207;
wire n_22208;
wire n_22209;
wire n_22210;
wire n_22211;
wire n_22212;
wire n_22213;
wire n_22214;
wire n_22215;
wire n_22216;
wire n_22217;
wire n_22218;
wire n_22219;
wire n_22220;
wire n_22221;
wire n_22222;
wire n_22223;
wire n_22224;
wire n_22225;
wire n_22226;
wire n_22227;
wire n_22228;
wire n_22229;
wire n_22230;
wire n_22231;
wire n_22232;
wire n_22233;
wire n_22234;
wire n_22235;
wire n_22236;
wire n_22237;
wire n_22238;
wire n_22239;
wire n_22240;
wire n_22241;
wire n_22242;
wire n_22243;
wire n_22244;
wire n_22245;
wire n_22246;
wire n_22247;
wire n_22248;
wire n_22249;
wire n_22250;
wire n_22251;
wire n_22252;
wire n_22253;
wire n_22254;
wire n_22255;
wire n_22256;
wire n_22257;
wire n_22258;
wire n_22259;
wire n_22260;
wire n_22261;
wire n_22262;
wire n_22263;
wire n_22264;
wire n_22265;
wire n_22266;
wire n_22267;
wire n_22268;
wire n_22269;
wire n_22270;
wire n_22271;
wire n_22272;
wire n_22273;
wire n_22274;
wire n_22275;
wire n_22276;
wire n_22277;
wire n_22278;
wire n_22279;
wire n_22280;
wire n_22281;
wire n_22282;
wire n_22283;
wire n_22284;
wire n_22285;
wire n_22286;
wire n_22287;
wire n_22288;
wire n_22289;
wire n_22290;
wire n_22291;
wire n_22292;
wire n_22293;
wire n_22294;
wire n_22295;
wire n_22296;
wire n_22297;
wire n_22298;
wire n_22299;
wire n_22300;
wire n_22301;
wire n_22302;
wire n_22303;
wire n_22304;
wire n_22305;
wire n_22306;
wire n_22307;
wire n_22308;
wire n_22309;
wire n_22310;
wire n_22311;
wire n_22312;
wire n_22313;
wire n_22314;
wire n_22315;
wire n_22316;
wire n_22317;
wire n_22318;
wire n_22319;
wire n_22320;
wire n_22321;
wire n_22322;
wire n_22323;
wire n_22324;
wire n_22325;
wire n_22326;
wire n_22327;
wire n_22328;
wire n_22329;
wire n_22330;
wire n_22331;
wire n_22332;
wire n_22333;
wire n_22334;
wire n_22335;
wire n_22336;
wire n_22337;
wire n_22338;
wire n_22339;
wire n_22340;
wire n_22341;
wire n_22342;
wire n_22343;
wire n_22344;
wire n_22345;
wire n_22346;
wire n_22347;
wire n_22348;
wire n_22349;
wire n_22350;
wire n_22351;
wire n_22352;
wire n_22353;
wire n_22354;
wire n_22355;
wire n_22356;
wire n_22357;
wire n_22358;
wire n_22359;
wire n_22360;
wire n_22361;
wire n_22362;
wire n_22363;
wire n_22364;
wire n_22365;
wire n_22366;
wire n_22367;
wire n_22368;
wire n_22369;
wire n_22370;
wire n_22371;
wire n_22372;
wire n_22373;
wire n_22374;
wire n_22375;
wire n_22376;
wire n_22377;
wire n_22378;
wire n_22379;
wire n_22380;
wire n_22381;
wire n_22382;
wire n_22383;
wire n_22384;
wire n_22385;
wire n_22386;
wire n_22387;
wire n_22388;
wire n_22389;
wire n_22390;
wire n_22391;
wire n_22392;
wire n_22393;
wire n_22394;
wire n_22395;
wire n_22396;
wire n_22397;
wire n_22398;
wire n_22399;
wire n_22400;
wire n_22401;
wire n_22402;
wire n_22403;
wire n_22404;
wire n_22405;
wire n_22406;
wire n_22407;
wire n_22408;
wire n_22409;
wire n_22410;
wire n_22411;
wire n_22412;
wire n_22413;
wire n_22414;
wire n_22415;
wire n_22416;
wire n_22417;
wire n_22418;
wire n_22419;
wire n_22420;
wire n_22421;
wire n_22422;
wire n_22423;
wire n_22424;
wire n_22425;
wire n_22426;
wire n_22427;
wire n_22428;
wire n_22429;
wire n_22430;
wire n_22431;
wire n_22432;
wire n_22433;
wire n_22434;
wire n_22435;
wire n_22436;
wire n_22437;
wire n_22438;
wire n_22439;
wire n_22440;
wire n_22441;
wire n_22442;
wire n_22443;
wire n_22444;
wire n_22445;
wire n_22446;
wire n_22447;
wire n_22448;
wire n_22449;
wire n_22450;
wire n_22451;
wire n_22452;
wire n_22453;
wire n_22454;
wire n_22455;
wire n_22456;
wire n_22457;
wire n_22458;
wire n_22459;
wire n_22460;
wire n_22461;
wire n_22462;
wire n_22463;
wire n_22464;
wire n_22465;
wire n_22466;
wire n_22467;
wire n_22468;
wire n_22469;
wire n_22470;
wire n_22471;
wire n_22472;
wire n_22473;
wire n_22474;
wire n_22475;
wire n_22476;
wire n_22477;
wire n_22478;
wire n_22479;
wire n_22480;
wire n_22481;
wire n_22482;
wire n_22483;
wire n_22484;
wire n_22485;
wire n_22486;
wire n_22487;
wire n_22488;
wire n_22489;
wire n_22490;
wire n_22491;
wire n_22492;
wire n_22493;
wire n_22494;
wire n_22495;
wire n_22496;
wire n_22497;
wire n_22498;
wire n_22499;
wire n_22500;
wire n_22501;
wire n_22502;
wire n_22503;
wire n_22504;
wire n_22505;
wire n_22506;
wire n_22507;
wire n_22508;
wire n_22509;
wire n_22510;
wire n_22511;
wire n_22512;
wire n_22513;
wire n_22514;
wire n_22515;
wire n_22516;
wire n_22517;
wire n_22518;
wire n_22519;
wire n_22520;
wire n_22521;
wire n_22522;
wire n_22523;
wire n_22524;
wire n_22525;
wire n_22526;
wire n_22527;
wire n_22528;
wire n_22529;
wire n_22530;
wire n_22531;
wire n_22532;
wire n_22533;
wire n_22534;
wire n_22535;
wire n_22536;
wire n_22537;
wire n_22538;
wire n_22539;
wire n_22540;
wire n_22541;
wire n_22542;
wire n_22543;
wire n_22544;
wire n_22545;
wire n_22546;
wire n_22547;
wire n_22548;
wire n_22549;
wire n_22550;
wire n_22551;
wire n_22552;
wire n_22553;
wire n_22554;
wire n_22555;
wire n_22556;
wire n_22557;
wire n_22558;
wire n_22559;
wire n_22560;
wire n_22561;
wire n_22562;
wire n_22563;
wire n_22564;
wire n_22565;
wire n_22566;
wire n_22567;
wire n_22568;
wire n_22569;
wire n_22570;
wire n_22571;
wire n_22572;
wire n_22573;
wire n_22574;
wire n_22575;
wire n_22576;
wire n_22577;
wire n_22578;
wire n_22579;
wire n_22580;
wire n_22581;
wire n_22582;
wire n_22583;
wire n_22584;
wire n_22585;
wire n_22586;
wire n_22587;
wire n_22588;
wire n_22589;
wire n_22590;
wire n_22591;
wire n_22592;
wire n_22593;
wire n_22594;
wire n_22595;
wire n_22596;
wire n_22597;
wire n_22598;
wire n_22599;
wire n_22600;
wire n_22601;
wire n_22602;
wire n_22603;
wire n_22604;
wire n_22605;
wire n_22606;
wire n_22607;
wire n_22608;
wire n_22609;
wire n_22610;
wire n_22611;
wire n_22612;
wire n_22613;
wire n_22614;
wire n_22615;
wire n_22616;
wire n_22617;
wire n_22618;
wire n_22619;
wire n_22620;
wire n_22621;
wire n_22622;
wire n_22623;
wire n_22624;
wire n_22625;
wire n_22626;
wire n_22627;
wire n_22628;
wire n_22629;
wire n_22630;
wire n_22631;
wire n_22632;
wire n_22633;
wire n_22634;
wire n_22635;
wire n_22636;
wire n_22637;
wire n_22638;
wire n_22639;
wire n_22640;
wire n_22641;
wire n_22642;
wire n_22643;
wire n_22644;
wire n_22645;
wire n_22646;
wire n_22647;
wire n_22648;
wire n_22649;
wire n_22650;
wire n_22651;
wire n_22652;
wire n_22653;
wire n_22654;
wire n_22655;
wire n_22656;
wire n_22657;
wire n_22658;
wire n_22659;
wire n_22660;
wire n_22661;
wire n_22662;
wire n_22663;
wire n_22664;
wire n_22665;
wire n_22666;
wire n_22667;
wire n_22668;
wire n_22669;
wire n_22670;
wire n_22671;
wire n_22672;
wire n_22673;
wire n_22674;
wire n_22675;
wire n_22676;
wire n_22677;
wire n_22678;
wire n_22679;
wire n_22680;
wire n_22681;
wire n_22682;
wire n_22683;
wire n_22684;
wire n_22685;
wire n_22686;
wire n_22687;
wire n_22688;
wire n_22689;
wire n_22690;
wire n_22691;
wire n_22692;
wire n_22693;
wire n_22694;
wire n_22695;
wire n_22696;
wire n_22697;
wire n_22698;
wire n_22699;
wire n_22700;
wire n_22701;
wire n_22702;
wire n_22703;
wire n_22704;
wire n_22705;
wire n_22706;
wire n_22707;
wire n_22708;
wire n_22709;
wire n_22710;
wire n_22711;
wire n_22712;
wire n_22713;
wire n_22714;
wire n_22715;
wire n_22716;
wire n_22717;
wire n_22718;
wire n_22719;
wire n_22720;
wire n_22721;
wire n_22722;
wire n_22723;
wire n_22724;
wire n_22725;
wire n_22726;
wire n_22727;
wire n_22728;
wire n_22729;
wire n_22730;
wire n_22731;
wire n_22732;
wire n_22733;
wire n_22734;
wire n_22735;
wire n_22736;
wire n_22737;
wire n_22738;
wire n_22739;
wire n_22740;
wire n_22741;
wire n_22742;
wire n_22743;
wire n_22744;
wire n_22745;
wire n_22746;
wire n_22747;
wire n_22748;
wire n_22749;
wire n_22750;
wire n_22751;
wire n_22752;
wire n_22753;
wire n_22754;
wire n_22755;
wire n_22756;
wire n_22757;
wire n_22758;
wire n_22759;
wire n_22760;
wire n_22761;
wire n_22762;
wire n_22763;
wire n_22764;
wire n_22765;
wire n_22766;
wire n_22767;
wire n_22768;
wire n_22769;
wire n_22770;
wire n_22771;
wire n_22772;
wire n_22773;
wire n_22774;
wire n_22775;
wire n_22776;
wire n_22777;
wire n_22778;
wire n_22779;
wire n_22780;
wire n_22781;
wire n_22782;
wire n_22783;
wire n_22784;
wire n_22785;
wire n_22786;
wire n_22787;
wire n_22788;
wire n_22789;
wire n_22790;
wire n_22791;
wire n_22792;
wire n_22793;
wire n_22794;
wire n_22795;
wire n_22796;
wire n_22797;
wire n_22798;
wire n_22799;
wire n_22800;
wire n_22801;
wire n_22802;
wire n_22803;
wire n_22804;
wire n_22805;
wire n_22806;
wire n_22807;
wire n_22808;
wire n_22809;
wire n_22810;
wire n_22811;
wire n_22812;
wire n_22813;
wire n_22814;
wire n_22815;
wire n_22816;
wire n_22817;
wire n_22818;
wire n_22819;
wire n_22820;
wire n_22821;
wire n_22822;
wire n_22823;
wire n_22824;
wire n_22825;
wire n_22826;
wire n_22827;
wire n_22828;
wire n_22829;
wire n_22830;
wire n_22831;
wire n_22832;
wire n_22833;
wire n_22834;
wire n_22835;
wire n_22836;
wire n_22837;
wire n_22838;
wire n_22839;
wire n_22840;
wire n_22841;
wire n_22842;
wire n_22843;
wire n_22844;
wire n_22845;
wire n_22846;
wire n_22847;
wire n_22848;
wire n_22849;
wire n_22850;
wire n_22851;
wire n_22852;
wire n_22853;
wire n_22854;
wire n_22855;
wire n_22856;
wire n_22857;
wire n_22858;
wire n_22859;
wire n_22860;
wire n_22861;
wire n_22862;
wire n_22863;
wire n_22864;
wire n_22865;
wire n_22866;
wire n_22867;
wire n_22868;
wire n_22869;
wire n_22870;
wire n_22871;
wire n_22872;
wire n_22873;
wire n_22874;
wire n_22875;
wire n_22876;
wire n_22877;
wire n_22878;
wire n_22879;
wire n_22880;
wire n_22881;
wire n_22882;
wire n_22883;
wire n_22884;
wire n_22885;
wire n_22886;
wire n_22887;
wire n_22888;
wire n_22889;
wire n_22890;
wire n_22891;
wire n_22892;
wire n_22893;
wire n_22894;
wire n_22895;
wire n_22896;
wire n_22897;
wire n_22898;
wire n_22899;
wire n_22900;
wire n_22901;
wire n_22902;
wire n_22903;
wire n_22904;
wire n_22905;
wire n_22906;
wire n_22907;
wire n_22908;
wire n_22909;
wire n_22910;
wire n_22911;
wire n_22912;
wire n_22913;
wire n_22914;
wire n_22915;
wire n_22916;
wire n_22917;
wire n_22918;
wire n_22919;
wire n_22920;
wire n_22921;
wire n_22922;
wire n_22923;
wire n_22924;
wire n_22925;
wire n_22926;
wire n_22927;
wire n_22928;
wire n_22929;
wire n_22930;
wire n_22931;
wire n_22932;
wire n_22933;
wire n_22934;
wire n_22935;
wire n_22936;
wire n_22937;
wire n_22938;
wire n_22939;
wire n_22940;
wire n_22941;
wire n_22942;
wire n_22943;
wire n_22944;
wire n_22945;
wire n_22946;
wire n_22947;
wire n_22948;
wire n_22949;
wire n_22950;
wire n_22951;
wire n_22952;
wire n_22953;
wire n_22954;
wire n_22955;
wire n_22956;
wire n_22957;
wire n_22958;
wire n_22959;
wire n_22960;
wire n_22961;
wire n_22962;
wire n_22963;
wire n_22964;
wire n_22965;
wire n_22966;
wire n_22967;
wire n_22968;
wire n_22969;
wire n_22970;
wire n_22971;
wire n_22972;
wire n_22973;
wire n_22974;
wire n_22975;
wire n_22976;
wire n_22977;
wire n_22978;
wire n_22979;
wire n_22980;
wire n_22981;
wire n_22982;
wire n_22983;
wire n_22984;
wire n_22985;
wire n_22986;
wire n_22987;
wire n_22988;
wire n_22989;
wire n_22990;
wire n_22991;
wire n_22992;
wire n_22993;
wire n_22994;
wire n_22995;
wire n_22996;
wire n_22997;
wire n_22998;
wire n_22999;
wire n_23000;
wire n_23001;
wire n_23002;
wire n_23003;
wire n_23004;
wire n_23005;
wire n_23006;
wire n_23007;
wire n_23008;
wire n_23009;
wire n_23010;
wire n_23011;
wire n_23012;
wire n_23013;
wire n_23014;
wire n_23015;
wire n_23016;
wire n_23017;
wire n_23018;
wire n_23019;
wire n_23020;
wire n_23021;
wire n_23022;
wire n_23023;
wire n_23024;
wire n_23025;
wire n_23026;
wire n_23027;
wire n_23028;
wire n_23029;
wire n_23030;
wire n_23031;
wire n_23032;
wire n_23033;
wire n_23034;
wire n_23035;
wire n_23036;
wire n_23037;
wire n_23038;
wire n_23039;
wire n_23040;
wire n_23041;
wire n_23042;
wire n_23043;
wire n_23044;
wire n_23045;
wire n_23046;
wire n_23047;
wire n_23048;
wire n_23049;
wire n_23050;
wire n_23051;
wire n_23052;
wire n_23053;
wire n_23054;
wire n_23055;
wire n_23056;
wire n_23057;
wire n_23058;
wire n_23059;
wire n_23060;
wire n_23061;
wire n_23062;
wire n_23063;
wire n_23064;
wire n_23065;
wire n_23066;
wire n_23067;
wire n_23068;
wire n_23069;
wire n_23070;
wire n_23071;
wire n_23072;
wire n_23073;
wire n_23074;
wire n_23075;
wire n_23076;
wire n_23077;
wire n_23078;
wire n_23079;
wire n_23080;
wire n_23081;
wire n_23082;
wire n_23083;
wire n_23084;
wire n_23085;
wire n_23086;
wire n_23087;
wire n_23088;
wire n_23089;
wire n_23090;
wire n_23091;
wire n_23092;
wire n_23093;
wire n_23094;
wire n_23095;
wire n_23096;
wire n_23097;
wire n_23098;
wire n_23099;
wire n_23100;
wire n_23101;
wire n_23102;
wire n_23103;
wire n_23104;
wire n_23105;
wire n_23106;
wire n_23107;
wire n_23108;
wire n_23109;
wire n_23110;
wire n_23111;
wire n_23112;
wire n_23113;
wire n_23114;
wire n_23115;
wire n_23116;
wire n_23117;
wire n_23118;
wire n_23119;
wire n_23120;
wire n_23121;
wire n_23122;
wire n_23123;
wire n_23124;
wire n_23125;
wire n_23126;
wire n_23127;
wire n_23128;
wire n_23129;
wire n_23130;
wire n_23131;
wire n_23132;
wire n_23133;
wire n_23134;
wire n_23135;
wire n_23136;
wire n_23137;
wire n_23138;
wire n_23139;
wire n_23140;
wire n_23141;
wire n_23142;
wire n_23143;
wire n_23144;
wire n_23145;
wire n_23146;
wire n_23147;
wire n_23148;
wire n_23149;
wire n_23150;
wire n_23151;
wire n_23152;
wire n_23153;
wire n_23154;
wire n_23155;
wire n_23156;
wire n_23157;
wire n_23158;
wire n_23159;
wire n_23160;
wire n_23161;
wire n_23162;
wire n_23163;
wire n_23164;
wire n_23165;
wire n_23166;
wire n_23167;
wire n_23168;
wire n_23169;
wire n_23170;
wire n_23171;
wire n_23172;
wire n_23173;
wire n_23174;
wire n_23175;
wire n_23176;
wire n_23177;
wire n_23178;
wire n_23179;
wire n_23180;
wire n_23181;
wire n_23182;
wire n_23183;
wire n_23184;
wire n_23185;
wire n_23186;
wire n_23187;
wire n_23188;
wire n_23189;
wire n_23190;
wire n_23191;
wire n_23192;
wire n_23193;
wire n_23194;
wire n_23195;
wire n_23196;
wire n_23197;
wire n_23198;
wire n_23199;
wire n_23200;
wire n_23201;
wire n_23202;
wire n_23203;
wire n_23204;
wire n_23205;
wire n_23206;
wire n_23207;
wire n_23208;
wire n_23209;
wire n_23210;
wire n_23211;
wire n_23212;
wire n_23213;
wire n_23214;
wire n_23215;
wire n_23216;
wire n_23217;
wire n_23218;
wire n_23219;
wire n_23220;
wire n_23221;
wire n_23222;
wire n_23223;
wire n_23224;
wire n_23225;
wire n_23226;
wire n_23227;
wire n_23228;
wire n_23229;
wire n_23230;
wire n_23231;
wire n_23232;
wire n_23233;
wire n_23234;
wire n_23235;
wire n_23236;
wire n_23237;
wire n_23238;
wire n_23239;
wire n_23240;
wire n_23241;
wire n_23242;
wire n_23243;
wire n_23244;
wire n_23245;
wire n_23246;
wire n_23247;
wire n_23248;
wire n_23249;
wire n_23250;
wire n_23251;
wire n_23252;
wire n_23253;
wire n_23254;
wire n_23255;
wire n_23256;
wire n_23257;
wire n_23258;
wire n_23259;
wire n_23260;
wire n_23261;
wire n_23262;
wire n_23263;
wire n_23264;
wire n_23265;
wire n_23266;
wire n_23267;
wire n_23268;
wire n_23269;
wire n_23270;
wire n_23271;
wire n_23272;
wire n_23273;
wire n_23274;
wire n_23275;
wire n_23276;
wire n_23277;
wire n_23278;
wire n_23279;
wire n_23280;
wire n_23281;
wire n_23282;
wire n_23283;
wire n_23284;
wire n_23285;
wire n_23286;
wire n_23287;
wire n_23288;
wire n_23289;
wire n_23290;
wire n_23291;
wire n_23292;
wire n_23293;
wire n_23294;
wire n_23295;
wire n_23296;
wire n_23297;
wire n_23298;
wire n_23299;
wire n_23300;
wire n_23301;
wire n_23302;
wire n_23303;
wire n_23304;
wire n_23305;
wire n_23306;
wire n_23307;
wire n_23308;
wire n_23309;
wire n_23310;
wire n_23311;
wire n_23312;
wire n_23313;
wire n_23314;
wire n_23315;
wire n_23316;
wire n_23317;
wire n_23318;
wire n_23319;
wire n_23320;
wire n_23321;
wire n_23322;
wire n_23323;
wire n_23324;
wire n_23325;
wire n_23326;
wire n_23327;
wire n_23328;
wire n_23329;
wire n_23330;
wire n_23331;
wire n_23332;
wire n_23333;
wire n_23334;
wire n_23335;
wire n_23336;
wire n_23337;
wire n_23338;
wire n_23339;
wire n_23340;
wire n_23341;
wire n_23342;
wire n_23343;
wire n_23344;
wire n_23345;
wire n_23346;
wire n_23347;
wire n_23348;
wire n_23349;
wire n_23350;
wire n_23351;
wire n_23352;
wire n_23353;
wire n_23354;
wire n_23355;
wire n_23356;
wire n_23357;
wire n_23358;
wire n_23359;
wire n_23360;
wire n_23361;
wire n_23362;
wire n_23363;
wire n_23364;
wire n_23365;
wire n_23366;
wire n_23367;
wire n_23368;
wire n_23369;
wire n_23370;
wire n_23371;
wire n_23372;
wire n_23373;
wire n_23374;
wire n_23375;
wire n_23376;
wire n_23377;
wire n_23378;
wire n_23379;
wire n_23380;
wire n_23381;
wire n_23382;
wire n_23383;
wire n_23384;
wire n_23385;
wire n_23386;
wire n_23387;
wire n_23388;
wire n_23389;
wire n_23390;
wire n_23391;
wire n_23392;
wire n_23393;
wire n_23394;
wire n_23395;
wire n_23396;
wire n_23397;
wire n_23398;
wire n_23399;
wire n_23400;
wire n_23401;
wire n_23402;
wire n_23403;
wire n_23404;
wire n_23405;
wire n_23406;
wire n_23407;
wire n_23408;
wire n_23409;
wire n_23410;
wire n_23411;
wire n_23412;
wire n_23413;
wire n_23414;
wire n_23415;
wire n_23416;
wire n_23417;
wire n_23418;
wire n_23419;
wire n_23420;
wire n_23421;
wire n_23422;
wire n_23423;
wire n_23424;
wire n_23425;
wire n_23426;
wire n_23427;
wire n_23428;
wire n_23429;
wire n_23430;
wire n_23431;
wire n_23432;
wire n_23433;
wire n_23434;
wire n_23435;
wire n_23436;
wire n_23437;
wire n_23438;
wire n_23439;
wire n_23440;
wire n_23441;
wire n_23442;
wire n_23443;
wire n_23444;
wire n_23445;
wire n_23446;
wire n_23447;
wire n_23448;
wire n_23449;
wire n_23450;
wire n_23451;
wire n_23452;
wire n_23453;
wire n_23454;
wire n_23455;
wire n_23456;
wire n_23457;
wire n_23458;
wire n_23459;
wire n_23460;
wire n_23461;
wire n_23462;
wire n_23463;
wire n_23464;
wire n_23465;
wire n_23466;
wire n_23467;
wire n_23468;
wire n_23469;
wire n_23470;
wire n_23471;
wire n_23472;
wire n_23473;
wire n_23474;
wire n_23475;
wire n_23476;
wire n_23477;
wire n_23478;
wire n_23479;
wire n_23480;
wire n_23481;
wire n_23482;
wire n_23483;
wire n_23484;
wire n_23485;
wire n_23486;
wire n_23487;
wire n_23488;
wire n_23489;
wire n_23490;
wire n_23491;
wire n_23492;
wire n_23493;
wire n_23494;
wire n_23495;
wire n_23496;
wire n_23497;
wire n_23498;
wire n_23499;
wire n_23500;
wire n_23501;
wire n_23502;
wire n_23503;
wire n_23504;
wire n_23505;
wire n_23506;
wire n_23507;
wire n_23508;
wire n_23509;
wire n_23510;
wire n_23511;
wire n_23512;
wire n_23513;
wire n_23514;
wire n_23515;
wire n_23516;
wire n_23517;
wire n_23518;
wire n_23519;
wire n_23520;
wire n_23521;
wire n_23522;
wire n_23523;
wire n_23524;
wire n_23525;
wire n_23526;
wire n_23527;
wire n_23528;
wire n_23529;
wire n_23530;
wire n_23531;
wire n_23532;
wire n_23533;
wire n_23534;
wire n_23535;
wire n_23536;
wire n_23537;
wire n_23538;
wire n_23539;
wire n_23540;
wire n_23541;
wire n_23542;
wire n_23543;
wire n_23544;
wire n_23545;
wire n_23546;
wire n_23547;
wire n_23548;
wire n_23549;
wire n_23550;
wire n_23551;
wire n_23552;
wire n_23553;
wire n_23554;
wire n_23555;
wire n_23556;
wire n_23557;
wire n_23558;
wire n_23559;
wire n_23560;
wire n_23561;
wire n_23562;
wire n_23563;
wire n_23564;
wire n_23565;
wire n_23566;
wire n_23567;
wire n_23568;
wire n_23569;
wire n_23570;
wire n_23571;
wire n_23572;
wire n_23573;
wire n_23574;
wire n_23575;
wire n_23576;
wire n_23577;
wire n_23578;
wire n_23579;
wire n_23580;
wire n_23581;
wire n_23582;
wire n_23583;
wire n_23584;
wire n_23585;
wire n_23586;
wire n_23587;
wire n_23588;
wire n_23589;
wire n_23590;
wire n_23591;
wire n_23592;
wire n_23593;
wire n_23594;
wire n_23595;
wire n_23596;
wire n_23597;
wire n_23598;
wire n_23599;
wire n_23600;
wire n_23601;
wire n_23602;
wire n_23603;
wire n_23604;
wire n_23605;
wire n_23606;
wire n_23607;
wire n_23608;
wire n_23609;
wire n_23610;
wire n_23611;
wire n_23612;
wire n_23613;
wire n_23614;
wire n_23615;
wire n_23616;
wire n_23617;
wire n_23618;
wire n_23619;
wire n_23620;
wire n_23621;
wire n_23622;
wire n_23623;
wire n_23624;
wire n_23625;
wire n_23626;
wire n_23627;
wire n_23628;
wire n_23629;
wire n_23630;
wire n_23631;
wire n_23632;
wire n_23633;
wire n_23634;
wire n_23635;
wire n_23636;
wire n_23637;
wire n_23638;
wire n_23639;
wire n_23640;
wire n_23641;
wire n_23642;
wire n_23643;
wire n_23644;
wire n_23645;
wire n_23646;
wire n_23647;
wire n_23648;
wire n_23649;
wire n_23650;
wire n_23651;
wire n_23652;
wire n_23653;
wire n_23654;
wire n_23655;
wire n_23656;
wire n_23657;
wire n_23658;
wire n_23659;
wire n_23660;
wire n_23661;
wire n_23662;
wire n_23663;
wire n_23664;
wire n_23665;
wire n_23666;
wire n_23667;
wire n_23668;
wire n_23669;
wire n_23670;
wire n_23671;
wire n_23672;
wire n_23673;
wire n_23674;
wire n_23675;
wire n_23676;
wire n_23677;
wire n_23678;
wire n_23679;
wire n_23680;
wire n_23681;
wire n_23682;
wire n_23683;
wire n_23684;
wire n_23685;
wire n_23686;
wire n_23687;
wire n_23688;
wire n_23689;
wire n_23690;
wire n_23691;
wire n_23692;
wire n_23693;
wire n_23694;
wire n_23695;
wire n_23696;
wire n_23697;
wire n_23698;
wire n_23699;
wire n_23700;
wire n_23701;
wire n_23702;
wire n_23703;
wire n_23704;
wire n_23705;
wire n_23706;
wire n_23707;
wire n_23708;
wire n_23709;
wire n_23710;
wire n_23711;
wire n_23712;
wire n_23713;
wire n_23714;
wire n_23715;
wire n_23716;
wire n_23717;
wire n_23718;
wire n_23719;
wire n_23720;
wire n_23721;
wire n_23722;
wire n_23723;
wire n_23724;
wire n_23725;
wire n_23726;
wire n_23727;
wire n_23728;
wire n_23729;
wire n_23730;
wire n_23731;
wire n_23732;
wire n_23733;
wire n_23734;
wire n_23735;
wire n_23736;
wire n_23737;
wire n_23738;
wire n_23739;
wire n_23740;
wire n_23741;
wire n_23742;
wire n_23743;
wire n_23744;
wire n_23745;
wire n_23746;
wire n_23747;
wire n_23748;
wire n_23749;
wire n_23750;
wire n_23751;
wire n_23752;
wire n_23753;
wire n_23754;
wire n_23755;
wire n_23756;
wire n_23757;
wire n_23758;
wire n_23759;
wire n_23760;
wire n_23761;
wire n_23762;
wire n_23763;
wire n_23764;
wire n_23765;
wire n_23766;
wire n_23767;
wire n_23768;
wire n_23769;
wire n_23770;
wire n_23771;
wire n_23772;
wire n_23773;
wire n_23774;
wire n_23775;
wire n_23776;
wire n_23777;
wire n_23778;
wire n_23779;
wire n_23780;
wire n_23781;
wire n_23782;
wire n_23783;
wire n_23784;
wire n_23785;
wire n_23786;
wire n_23787;
wire n_23788;
wire n_23789;
wire n_23790;
wire n_23791;
wire n_23792;
wire n_23793;
wire n_23794;
wire n_23795;
wire n_23796;
wire n_23797;
wire n_23798;
wire n_23799;
wire n_23800;
wire n_23801;
wire n_23802;
wire n_23803;
wire n_23804;
wire n_23805;
wire n_23806;
wire n_23807;
wire n_23808;
wire n_23809;
wire n_23810;
wire n_23811;
wire n_23812;
wire n_23813;
wire n_23814;
wire n_23815;
wire n_23816;
wire n_23817;
wire n_23818;
wire n_23819;
wire n_23820;
wire n_23821;
wire n_23822;
wire n_23823;
wire n_23824;
wire n_23825;
wire n_23826;
wire n_23827;
wire n_23828;
wire n_23829;
wire n_23830;
wire n_23831;
wire n_23832;
wire n_23833;
wire n_23834;
wire n_23835;
wire n_23836;
wire n_23837;
wire n_23838;
wire n_23839;
wire n_23840;
wire n_23841;
wire n_23842;
wire n_23843;
wire n_23844;
wire n_23845;
wire n_23846;
wire n_23847;
wire n_23848;
wire n_23849;
wire n_23850;
wire n_23851;
wire n_23852;
wire n_23853;
wire n_23854;
wire n_23855;
wire n_23856;
wire n_23857;
wire n_23858;
wire n_23859;
wire n_23860;
wire n_23861;
wire n_23862;
wire n_23863;
wire n_23864;
wire n_23865;
wire n_23866;
wire n_23867;
wire n_23868;
wire n_23869;
wire n_23870;
wire n_23871;
wire n_23872;
wire n_23873;
wire n_23874;
wire n_23875;
wire n_23876;
wire n_23877;
wire n_23878;
wire n_23879;
wire n_23880;
wire n_23881;
wire n_23882;
wire n_23883;
wire n_23884;
wire n_23885;
wire n_23886;
wire n_23887;
wire n_23888;
wire n_23889;
wire n_23890;
wire n_23891;
wire n_23892;
wire n_23893;
wire n_23894;
wire n_23895;
wire n_23896;
wire n_23897;
wire n_23898;
wire n_23899;
wire n_23900;
wire n_23901;
wire n_23902;
wire n_23903;
wire n_23904;
wire n_23905;
wire n_23906;
wire n_23907;
wire n_23908;
wire n_23909;
wire n_23910;
wire n_23911;
wire n_23912;
wire n_23913;
wire n_23914;
wire n_23915;
wire n_23916;
wire n_23917;
wire n_23918;
wire n_23919;
wire n_23920;
wire n_23921;
wire n_23922;
wire n_23923;
wire n_23924;
wire n_23925;
wire n_23926;
wire n_23927;
wire n_23928;
wire n_23929;
wire n_23930;
wire n_23931;
wire n_23932;
wire n_23933;
wire n_23934;
wire n_23935;
wire n_23936;
wire n_23937;
wire n_23938;
wire n_23939;
wire n_23940;
wire n_23941;
wire n_23942;
wire n_23943;
wire n_23944;
wire n_23945;
wire n_23946;
wire n_23947;
wire n_23948;
wire n_23949;
wire n_23950;
wire n_23951;
wire n_23952;
wire n_23953;
wire n_23954;
wire n_23955;
wire n_23956;
wire n_23957;
wire n_23958;
wire n_23959;
wire n_23960;
wire n_23961;
wire n_23962;
wire n_23963;
wire n_23964;
wire n_23965;
wire n_23966;
wire n_23967;
wire n_23968;
wire n_23969;
wire n_23970;
wire n_23971;
wire n_23972;
wire n_23973;
wire n_23974;
wire n_23975;
wire n_23976;
wire n_23977;
wire n_23978;
wire n_23979;
wire n_23980;
wire n_23981;
wire n_23982;
wire n_23983;
wire n_23984;
wire n_23985;
wire n_23986;
wire n_23987;
wire n_23988;
wire n_23989;
wire n_23990;
wire n_23991;
wire n_23992;
wire n_23993;
wire n_23994;
wire n_23995;
wire n_23996;
wire n_23997;
wire n_23998;
wire n_23999;
wire n_24000;
wire n_24001;
wire n_24002;
wire n_24003;
wire n_24004;
wire n_24005;
wire n_24006;
wire n_24007;
wire n_24008;
wire n_24009;
wire n_24010;
wire n_24011;
wire n_24012;
wire n_24013;
wire n_24014;
wire n_24015;
wire n_24016;
wire n_24017;
wire n_24018;
wire n_24019;
wire n_24020;
wire n_24021;
wire n_24022;
wire n_24023;
wire n_24024;
wire n_24025;
wire n_24026;
wire n_24027;
wire n_24028;
wire n_24029;
wire n_24030;
wire n_24031;
wire n_24032;
wire n_24033;
wire n_24034;
wire n_24035;
wire n_24036;
wire n_24037;
wire n_24038;
wire n_24039;
wire n_24040;
wire n_24041;
wire n_24042;
wire n_24043;
wire n_24044;
wire n_24045;
wire n_24046;
wire n_24047;
wire n_24048;
wire n_24049;
wire n_24050;
wire n_24051;
wire n_24052;
wire n_24053;
wire n_24054;
wire n_24055;
wire n_24056;
wire n_24057;
wire n_24058;
wire n_24059;
wire n_24060;
wire n_24061;
wire n_24062;
wire n_24063;
wire n_24064;
wire n_24065;
wire n_24066;
wire n_24067;
wire n_24068;
wire n_24069;
wire n_24070;
wire n_24071;
wire n_24072;
wire n_24073;
wire n_24074;
wire n_24075;
wire n_24076;
wire n_24077;
wire n_24078;
wire n_24079;
wire n_24080;
wire n_24081;
wire n_24082;
wire n_24083;
wire n_24084;
wire n_24085;
wire n_24086;
wire n_24087;
wire n_24088;
wire n_24089;
wire n_24090;
wire n_24091;
wire n_24092;
wire n_24093;
wire n_24094;
wire n_24095;
wire n_24096;
wire n_24097;
wire n_24098;
wire n_24099;
wire n_24100;
wire n_24101;
wire n_24102;
wire n_24103;
wire n_24104;
wire n_24105;
wire n_24106;
wire n_24107;
wire n_24108;
wire n_24109;
wire n_24110;
wire n_24111;
wire n_24112;
wire n_24113;
wire n_24114;
wire n_24115;
wire n_24116;
wire n_24117;
wire n_24118;
wire n_24119;
wire n_24120;
wire n_24121;
wire n_24122;
wire n_24123;
wire n_24124;
wire n_24125;
wire n_24126;
wire n_24127;
wire n_24128;
wire n_24129;
wire n_24130;
wire n_24131;
wire n_24132;
wire n_24133;
wire n_24134;
wire n_24135;
wire n_24136;
wire n_24137;
wire n_24138;
wire n_24139;
wire n_24140;
wire n_24141;
wire n_24142;
wire n_24143;
wire n_24144;
wire n_24145;
wire n_24146;
wire n_24147;
wire n_24148;
wire n_24149;
wire n_24150;
wire n_24151;
wire n_24152;
wire n_24153;
wire n_24154;
wire n_24155;
wire n_24156;
wire n_24157;
wire n_24158;
wire n_24159;
wire n_24160;
wire n_24161;
wire n_24162;
wire n_24163;
wire n_24164;
wire n_24165;
wire n_24166;
wire n_24167;
wire n_24168;
wire n_24169;
wire n_24170;
wire n_24171;
wire n_24172;
wire n_24173;
wire n_24174;
wire n_24175;
wire n_24176;
wire n_24177;
wire n_24178;
wire n_24179;
wire n_24180;
wire n_24181;
wire n_24182;
wire n_24183;
wire n_24184;
wire n_24185;
wire n_24186;
wire n_24187;
wire n_24188;
wire n_24189;
wire n_24190;
wire n_24191;
wire n_24192;
wire n_24193;
wire n_24194;
wire n_24195;
wire n_24196;
wire n_24197;
wire n_24198;
wire n_24199;
wire n_24200;
wire n_24201;
wire n_24202;
wire n_24203;
wire n_24204;
wire n_24205;
wire n_24206;
wire n_24207;
wire n_24208;
wire n_24209;
wire n_24210;
wire n_24211;
wire n_24212;
wire n_24213;
wire n_24214;
wire n_24215;
wire n_24216;
wire n_24217;
wire n_24218;
wire n_24219;
wire n_24220;
wire n_24221;
wire n_24222;
wire n_24223;
wire n_24224;
wire n_24225;
wire n_24226;
wire n_24227;
wire n_24228;
wire n_24229;
wire n_24230;
wire n_24231;
wire n_24232;
wire n_24233;
wire n_24234;
wire n_24235;
wire n_24236;
wire n_24237;
wire n_24238;
wire n_24239;
wire n_24240;
wire n_24241;
wire n_24242;
wire n_24243;
wire n_24244;
wire n_24245;
wire n_24246;
wire n_24247;
wire n_24248;
wire n_24249;
wire n_24250;
wire n_24251;
wire n_24252;
wire n_24253;
wire n_24254;
wire n_24255;
wire n_24256;
wire n_24257;
wire n_24258;
wire n_24259;
wire n_24260;
wire n_24261;
wire n_24262;
wire n_24263;
wire n_24264;
wire n_24265;
wire n_24266;
wire n_24267;
wire n_24268;
wire n_24269;
wire n_24270;
wire n_24271;
wire n_24272;
wire n_24273;
wire n_24274;
wire n_24275;
wire n_24276;
wire n_24277;
wire n_24278;
wire n_24279;
wire n_24280;
wire n_24281;
wire n_24282;
wire n_24283;
wire n_24284;
wire n_24285;
wire n_24286;
wire n_24287;
wire n_24288;
wire n_24289;
wire n_24290;
wire n_24291;
wire n_24292;
wire n_24293;
wire n_24294;
wire n_24295;
wire n_24296;
wire n_24297;
wire n_24298;
wire n_24299;
wire n_24300;
wire n_24301;
wire n_24302;
wire n_24303;
wire n_24304;
wire n_24305;
wire n_24306;
wire n_24307;
wire n_24308;
wire n_24309;
wire n_24310;
wire n_24311;
wire n_24312;
wire n_24313;
wire n_24314;
wire n_24315;
wire n_24316;
wire n_24317;
wire n_24318;
wire n_24319;
wire n_24320;
wire n_24321;
wire n_24322;
wire n_24323;
wire n_24324;
wire n_24325;
wire n_24326;
wire n_24327;
wire n_24328;
wire n_24329;
wire n_24330;
wire n_24331;
wire n_24332;
wire n_24333;
wire n_24334;
wire n_24335;
wire n_24336;
wire n_24337;
wire n_24338;
wire n_24339;
wire n_24340;
wire n_24341;
wire n_24342;
wire n_24343;
wire n_24344;
wire n_24345;
wire n_24346;
wire n_24347;
wire n_24348;
wire n_24349;
wire n_24350;
wire n_24351;
wire n_24352;
wire n_24353;
wire n_24354;
wire n_24355;
wire n_24356;
wire n_24357;
wire n_24358;
wire n_24359;
wire n_24360;
wire n_24361;
wire n_24362;
wire n_24363;
wire n_24364;
wire n_24365;
wire n_24366;
wire n_24367;
wire n_24368;
wire n_24369;
wire n_24370;
wire n_24371;
wire n_24372;
wire n_24373;
wire n_24374;
wire n_24375;
wire n_24376;
wire n_24377;
wire n_24378;
wire n_24379;
wire n_24380;
wire n_24381;
wire n_24382;
wire n_24383;
wire n_24384;
wire n_24385;
wire n_24386;
wire n_24387;
wire n_24388;
wire n_24389;
wire n_24390;
wire n_24391;
wire n_24392;
wire n_24393;
wire n_24394;
wire n_24395;
wire n_24396;
wire n_24397;
wire n_24398;
wire n_24399;
wire n_24400;
wire n_24401;
wire n_24402;
wire n_24403;
wire n_24404;
wire n_24405;
wire n_24406;
wire n_24407;
wire n_24408;
wire n_24409;
wire n_24410;
wire n_24411;
wire n_24412;
wire n_24413;
wire n_24414;
wire n_24415;
wire n_24416;
wire n_24417;
wire n_24418;
wire n_24419;
wire n_24420;
wire n_24421;
wire n_24422;
wire n_24423;
wire n_24424;
wire n_24425;
wire n_24426;
wire n_24427;
wire n_24428;
wire n_24429;
wire n_24430;
wire n_24431;
wire n_24432;
wire n_24433;
wire n_24434;
wire n_24435;
wire n_24436;
wire n_24437;
wire n_24438;
wire n_24439;
wire n_24440;
wire n_24441;
wire n_24442;
wire n_24443;
wire n_24444;
wire n_24445;
wire n_24446;
wire n_24447;
wire n_24448;
wire n_24449;
wire n_24450;
wire n_24451;
wire n_24452;
wire n_24453;
wire n_24454;
wire n_24455;
wire n_24456;
wire n_24457;
wire n_24458;
wire n_24459;
wire n_24460;
wire n_24461;
wire n_24462;
wire n_24463;
wire n_24464;
wire n_24465;
wire n_24466;
wire n_24467;
wire n_24468;
wire n_24469;
wire n_24470;
wire n_24471;
wire n_24472;
wire n_24473;
wire n_24474;
wire n_24475;
wire n_24476;
wire n_24477;
wire n_24478;
wire n_24479;
wire n_24480;
wire n_24481;
wire n_24482;
wire n_24483;
wire n_24484;
wire n_24485;
wire n_24486;
wire n_24487;
wire n_24488;
wire n_24489;
wire n_24490;
wire n_24491;
wire n_24492;
wire n_24493;
wire n_24494;
wire n_24495;
wire n_24496;
wire n_24497;
wire n_24498;
wire n_24499;
wire n_24500;
wire n_24501;
wire n_24502;
wire n_24503;
wire n_24504;
wire n_24505;
wire n_24506;
wire n_24507;
wire n_24508;
wire n_24509;
wire n_24510;
wire n_24511;
wire n_24512;
wire n_24513;
wire n_24514;
wire n_24515;
wire n_24516;
wire n_24517;
wire n_24518;
wire n_24519;
wire n_24520;
wire n_24521;
wire n_24522;
wire n_24523;
wire n_24524;
wire n_24525;
wire n_24526;
wire n_24527;
wire n_24528;
wire n_24529;
wire n_24530;
wire n_24531;
wire n_24532;
wire n_24533;
wire n_24534;
wire n_24535;
wire n_24536;
wire n_24537;
wire n_24538;
wire n_24539;
wire n_24540;
wire n_24541;
wire n_24542;
wire n_24543;
wire n_24544;
wire n_24545;
wire n_24546;
wire n_24547;
wire n_24548;
wire n_24549;
wire n_24550;
wire n_24551;
wire n_24552;
wire n_24553;
wire n_24554;
wire n_24555;
wire n_24556;
wire n_24557;
wire n_24558;
wire n_24559;
wire n_24560;
wire n_24561;
wire n_24562;
wire n_24563;
wire n_24564;
wire n_24565;
wire n_24566;
wire n_24567;
wire n_24568;
wire n_24569;
wire n_24570;
wire n_24571;
wire n_24572;
wire n_24573;
wire n_24574;
wire n_24575;
wire n_24576;
wire n_24577;
wire n_24578;
wire n_24579;
wire n_24580;
wire n_24581;
wire n_24582;
wire n_24583;
wire n_24584;
wire n_24585;
wire n_24586;
wire n_24587;
wire n_24588;
wire n_24589;
wire n_24590;
wire n_24591;
wire n_24592;
wire n_24593;
wire n_24594;
wire n_24595;
wire n_24596;
wire n_24597;
wire n_24598;
wire n_24599;
wire n_24600;
wire n_24601;
wire n_24602;
wire n_24603;
wire n_24604;
wire n_24605;
wire n_24606;
wire n_24607;
wire n_24608;
wire n_24609;
wire n_24610;
wire n_24611;
wire n_24612;
wire n_24613;
wire n_24614;
wire n_24615;
wire n_24616;
wire n_24617;
wire n_24618;
wire n_24619;
wire n_24620;
wire n_24621;
wire n_24622;
wire n_24623;
wire n_24624;
wire n_24625;
wire n_24626;
wire n_24627;
wire n_24628;
wire n_24629;
wire n_24630;
wire n_24631;
wire n_24632;
wire n_24633;
wire n_24634;
wire n_24635;
wire n_24636;
wire n_24637;
wire n_24638;
wire n_24639;
wire n_24640;
wire n_24641;
wire n_24642;
wire n_24643;
wire n_24644;
wire n_24645;
wire n_24646;
wire n_24647;
wire n_24648;
wire n_24649;
wire n_24650;
wire n_24651;
wire n_24652;
wire n_24653;
wire n_24654;
wire n_24655;
wire n_24656;
wire n_24657;
wire n_24658;
wire n_24659;
wire n_24660;
wire n_24661;
wire n_24662;
wire n_24663;
wire n_24664;
wire n_24665;
wire n_24666;
wire n_24667;
wire n_24668;
wire n_24669;
wire n_24670;
wire n_24671;
wire n_24672;
wire n_24673;
wire n_24674;
wire n_24675;
wire n_24676;
wire n_24677;
wire n_24678;
wire n_24679;
wire n_24680;
wire n_24681;
wire n_24682;
wire n_24683;
wire n_24684;
wire n_24685;
wire n_24686;
wire n_24687;
wire n_24688;
wire n_24689;
wire n_24690;
wire n_24691;
wire n_24692;
wire n_24693;
wire n_24694;
wire n_24695;
wire n_24696;
wire n_24697;
wire n_24698;
wire n_24699;
wire n_24700;
wire n_24701;
wire n_24702;
wire n_24703;
wire n_24704;
wire n_24705;
wire n_24706;
wire n_24707;
wire n_24708;
wire n_24709;
wire n_24710;
wire n_24711;
wire n_24712;
wire n_24713;
wire n_24714;
wire n_24715;
wire n_24716;
wire n_24717;
wire n_24718;
wire n_24719;
wire n_24720;
wire n_24721;
wire n_24722;
wire n_24723;
wire n_24724;
wire n_24725;
wire n_24726;
wire n_24727;
wire n_24728;
wire n_24729;
wire n_24730;
wire n_24731;
wire n_24732;
wire n_24733;
wire n_24734;
wire n_24735;
wire n_24736;
wire n_24737;
wire n_24738;
wire n_24739;
wire n_24740;
wire n_24741;
wire n_24742;
wire n_24743;
wire n_24744;
wire n_24745;
wire n_24746;
wire n_24747;
wire n_24748;
wire n_24749;
wire n_24750;
wire n_24751;
wire n_24752;
wire n_24753;
wire n_24754;
wire n_24755;
wire n_24756;
wire n_24757;
wire n_24758;
wire n_24759;
wire n_24760;
wire n_24761;
wire n_24762;
wire n_24763;
wire n_24764;
wire n_24765;
wire n_24766;
wire n_24767;
wire n_24768;
wire n_24769;
wire n_24770;
wire n_24771;
wire n_24772;
wire n_24773;
wire n_24774;
wire n_24775;
wire n_24776;
wire n_24777;
wire n_24778;
wire n_24779;
wire n_24780;
wire n_24781;
wire n_24782;
wire n_24783;
wire n_24784;
wire n_24785;
wire n_24786;
wire n_24787;
wire n_24788;
wire n_24789;
wire n_24790;
wire n_24791;
wire n_24792;
wire n_24793;
wire n_24794;
wire n_24795;
wire n_24796;
wire n_24797;
wire n_24798;
wire n_24799;
wire n_24800;
wire n_24801;
wire n_24802;
wire n_24803;
wire n_24804;
wire n_24805;
wire n_24806;
wire n_24807;
wire n_24808;
wire n_24809;
wire n_24810;
wire n_24811;
wire n_24812;
wire n_24813;
wire n_24814;
wire n_24815;
wire n_24816;
wire n_24817;
wire n_24818;
wire n_24819;
wire n_24820;
wire n_24821;
wire n_24822;
wire n_24823;
wire n_24824;
wire n_24825;
wire n_24826;
wire n_24827;
wire n_24828;
wire n_24829;
wire n_24830;
wire n_24831;
wire n_24832;
wire n_24833;
wire n_24834;
wire n_24835;
wire n_24836;
wire n_24837;
wire n_24838;
wire n_24839;
wire n_24840;
wire n_24841;
wire n_24842;
wire n_24843;
wire n_24844;
wire n_24845;
wire n_24846;
wire n_24847;
wire n_24848;
wire n_24849;
wire n_24850;
wire n_24851;
wire n_24852;
wire n_24853;
wire n_24854;
wire n_24855;
wire n_24856;
wire n_24857;
wire n_24858;
wire n_24859;
wire n_24860;
wire n_24861;
wire n_24862;
wire n_24863;
wire n_24864;
wire n_24865;
wire n_24866;
wire n_24867;
wire n_24868;
wire n_24869;
wire n_24870;
wire n_24871;
wire n_24872;
wire n_24873;
wire n_24874;
wire n_24875;
wire n_24876;
wire n_24877;
wire n_24878;
wire n_24879;
wire n_24880;
wire n_24881;
wire n_24882;
wire n_24883;
wire n_24884;
wire n_24885;
wire n_24886;
wire n_24887;
wire n_24888;
wire n_24889;
wire n_24890;
wire n_24891;
wire n_24892;
wire n_24893;
wire n_24894;
wire n_24895;
wire n_24896;
wire n_24897;
wire n_24898;
wire n_24899;
wire n_24900;
wire n_24901;
wire n_24902;
wire n_24903;
wire n_24904;
wire n_24905;
wire n_24906;
wire n_24907;
wire n_24908;
wire n_24909;
wire n_24910;
wire n_24911;
wire n_24912;
wire n_24913;
wire n_24914;
wire n_24915;
wire n_24916;
wire n_24917;
wire n_24918;
wire n_24919;
wire n_24920;
wire n_24921;
wire n_24922;
wire n_24923;
wire n_24924;
wire n_24925;
wire n_24926;
wire n_24927;
wire n_24928;
wire n_24929;
wire n_24930;
wire n_24931;
wire n_24932;
wire n_24933;
wire n_24934;
wire n_24935;
wire n_24936;
wire n_24937;
wire n_24938;
wire n_24939;
wire n_24940;
wire n_24941;
wire n_24942;
wire n_24943;
wire n_24944;
wire n_24945;
wire n_24946;
wire n_24947;
wire n_24948;
wire n_24949;
wire n_24950;
wire n_24951;
wire n_24952;
wire n_24953;
wire n_24954;
wire n_24955;
wire n_24956;
wire n_24957;
wire n_24958;
wire n_24959;
wire n_24960;
wire n_24961;
wire n_24962;
wire n_24963;
wire n_24964;
wire n_24965;
wire n_24966;
wire n_24967;
wire n_24968;
wire n_24969;
wire n_24970;
wire n_24971;
wire n_24972;
wire n_24973;
wire n_24974;
wire n_24975;
wire n_24976;
wire n_24977;
wire n_24978;
wire n_24979;
wire n_24980;
wire n_24981;
wire n_24982;
wire n_24983;
wire n_24984;
wire n_24985;
wire n_24986;
wire n_24987;
wire n_24988;
wire n_24989;
wire n_24990;
wire n_24991;
wire n_24992;
wire n_24993;
wire n_24994;
wire n_24995;
wire n_24996;
wire n_24997;
wire n_24998;
wire n_24999;
wire n_25000;
wire n_25001;
wire n_25002;
wire n_25003;
wire n_25004;
wire n_25005;
wire n_25006;
wire n_25007;
wire n_25008;
wire n_25009;
wire n_25010;
wire n_25011;
wire n_25012;
wire n_25013;
wire n_25014;
wire n_25015;
wire n_25016;
wire n_25017;
wire n_25018;
wire n_25019;
wire n_25020;
wire n_25021;
wire n_25022;
wire n_25023;
wire n_25024;
wire n_25025;
wire n_25026;
wire n_25027;
wire n_25028;
wire n_25029;
wire n_25030;
wire n_25031;
wire n_25032;
wire n_25033;
wire n_25034;
wire n_25035;
wire n_25036;
wire n_25037;
wire n_25038;
wire n_25039;
wire n_25040;
wire n_25041;
wire n_25042;
wire n_25043;
wire n_25044;
wire n_25045;
wire n_25046;
wire n_25047;
wire n_25048;
wire n_25049;
wire n_25050;
wire n_25051;
wire n_25052;
wire n_25053;
wire n_25054;
wire n_25055;
wire n_25056;
wire n_25057;
wire n_25058;
wire n_25059;
wire n_25060;
wire n_25061;
wire n_25062;
wire n_25063;
wire n_25064;
wire n_25065;
wire n_25066;
wire n_25067;
wire n_25068;
wire n_25069;
wire n_25070;
wire n_25071;
wire n_25072;
wire n_25073;
wire n_25074;
wire n_25075;
wire n_25076;
wire n_25077;
wire n_25078;
wire n_25079;
wire n_25080;
wire n_25081;
wire n_25082;
wire n_25083;
wire n_25084;
wire n_25085;
wire n_25086;
wire n_25087;
wire n_25088;
wire n_25089;
wire n_25090;
wire n_25091;
wire n_25092;
wire n_25093;
wire n_25094;
wire n_25095;
wire n_25096;
wire n_25097;
wire n_25098;
wire n_25099;
wire n_25100;
wire n_25101;
wire n_25102;
wire n_25103;
wire n_25104;
wire n_25105;
wire n_25106;
wire n_25107;
wire n_25108;
wire n_25109;
wire n_25110;
wire n_25111;
wire n_25112;
wire n_25113;
wire n_25114;
wire n_25115;
wire n_25116;
wire n_25117;
wire n_25118;
wire n_25119;
wire n_25120;
wire n_25121;
wire n_25122;
wire n_25123;
wire n_25124;
wire n_25125;
wire n_25126;
wire n_25127;
wire n_25128;
wire n_25129;
wire n_25130;
wire n_25131;
wire n_25132;
wire n_25133;
wire n_25134;
wire n_25135;
wire n_25136;
wire n_25137;
wire n_25138;
wire n_25139;
wire n_25140;
wire n_25141;
wire n_25142;
wire n_25143;
wire n_25144;
wire n_25145;
wire n_25146;
wire n_25147;
wire n_25148;
wire n_25149;
wire n_25150;
wire n_25151;
wire n_25152;
wire n_25153;
wire n_25154;
wire n_25155;
wire n_25156;
wire n_25157;
wire n_25158;
wire n_25159;
wire n_25160;
wire n_25161;
wire n_25162;
wire n_25163;
wire n_25164;
wire n_25165;
wire n_25166;
wire n_25167;
wire n_25168;
wire n_25169;
wire n_25170;
wire n_25171;
wire n_25172;
wire n_25173;
wire n_25174;
wire n_25175;
wire n_25176;
wire n_25177;
wire n_25178;
wire n_25179;
wire n_25180;
wire n_25181;
wire n_25182;
wire n_25183;
wire n_25184;
wire n_25185;
wire n_25186;
wire n_25187;
wire n_25188;
wire n_25189;
wire n_25190;
wire n_25191;
wire n_25192;
wire n_25193;
wire n_25194;
wire n_25195;
wire n_25196;
wire n_25197;
wire n_25198;
wire n_25199;
wire n_25200;
wire n_25201;
wire n_25202;
wire n_25203;
wire n_25204;
wire n_25205;
wire n_25206;
wire n_25207;
wire n_25208;
wire n_25209;
wire n_25210;
wire n_25211;
wire n_25212;
wire n_25213;
wire n_25214;
wire n_25215;
wire n_25216;
wire n_25217;
wire n_25218;
wire n_25219;
wire n_25220;
wire n_25221;
wire n_25222;
wire n_25223;
wire n_25224;
wire n_25225;
wire n_25226;
wire n_25227;
wire n_25228;
wire n_25229;
wire n_25230;
wire n_25231;
wire n_25232;
wire n_25233;
wire n_25234;
wire n_25235;
wire n_25236;
wire n_25237;
wire n_25238;
wire n_25239;
wire n_25240;
wire n_25241;
wire n_25242;
wire n_25243;
wire n_25244;
wire n_25245;
wire n_25246;
wire n_25247;
wire n_25248;
wire n_25249;
wire n_25250;
wire n_25251;
wire n_25252;
wire n_25253;
wire n_25254;
wire n_25255;
wire n_25256;
wire n_25257;
wire n_25258;
wire n_25259;
wire n_25260;
wire n_25261;
wire n_25262;
wire n_25263;
wire n_25264;
wire n_25265;
wire n_25266;
wire n_25267;
wire n_25268;
wire n_25269;
wire n_25270;
wire n_25271;
wire n_25272;
wire n_25273;
wire n_25274;
wire n_25275;
wire n_25276;
wire n_25277;
wire n_25278;
wire n_25279;
wire n_25280;
wire n_25281;
wire n_25282;
wire n_25283;
wire n_25284;
wire n_25285;
wire n_25286;
wire n_25287;
wire n_25288;
wire n_25289;
wire n_25290;
wire n_25291;
wire n_25292;
wire n_25293;
wire n_25294;
wire n_25295;
wire n_25296;
wire n_25297;
wire n_25298;
wire n_25299;
wire n_25300;
wire n_25301;
wire n_25302;
wire n_25303;
wire n_25304;
wire n_25305;
wire n_25306;
wire n_25307;
wire n_25308;
wire n_25309;
wire n_25310;
wire n_25311;
wire n_25312;
wire n_25313;
wire n_25314;
wire n_25315;
wire n_25316;
wire n_25317;
wire n_25318;
wire n_25319;
wire n_25320;
wire n_25321;
wire n_25322;
wire n_25323;
wire n_25324;
wire n_25325;
wire n_25326;
wire n_25327;
wire n_25328;
wire n_25329;
wire n_25330;
wire n_25331;
wire n_25332;
wire n_25333;
wire n_25334;
wire n_25335;
wire n_25336;
wire n_25337;
wire n_25338;
wire n_25339;
wire n_25340;
wire n_25341;
wire n_25342;
wire n_25343;
wire n_25344;
wire n_25345;
wire n_25346;
wire n_25347;
wire n_25348;
wire n_25349;
wire n_25350;
wire n_25351;
wire n_25352;
wire n_25353;
wire n_25354;
wire n_25355;
wire n_25356;
wire n_25357;
wire n_25358;
wire n_25359;
wire n_25360;
wire n_25361;
wire n_25362;
wire n_25363;
wire n_25364;
wire n_25365;
wire n_25366;
wire n_25367;
wire n_25368;
wire n_25369;
wire n_25370;
wire n_25371;
wire n_25372;
wire n_25373;
wire n_25374;
wire n_25375;
wire n_25376;
wire n_25377;
wire n_25378;
wire n_25379;
wire n_25380;
wire n_25381;
wire n_25382;
wire n_25383;
wire n_25384;
wire n_25385;
wire n_25386;
wire n_25387;
wire n_25388;
wire n_25389;
wire n_25390;
wire n_25391;
wire n_25392;
wire n_25393;
wire n_25394;
wire n_25395;
wire n_25396;
wire n_25397;
wire n_25398;
wire n_25399;
wire n_25400;
wire n_25401;
wire n_25402;
wire n_25403;
wire n_25404;
wire n_25405;
wire n_25406;
wire n_25407;
wire n_25408;
wire n_25409;
wire n_25410;
wire n_25411;
wire n_25412;
wire n_25413;
wire n_25414;
wire n_25415;
wire n_25416;
wire n_25417;
wire n_25418;
wire n_25419;
wire n_25420;
wire n_25421;
wire n_25422;
wire n_25423;
wire n_25424;
wire n_25425;
wire n_25426;
wire n_25427;
wire n_25428;
wire n_25429;
wire n_25430;
wire n_25431;
wire n_25432;
wire n_25433;
wire n_25434;
wire n_25435;
wire n_25436;
wire n_25437;
wire n_25438;
wire n_25439;
wire n_25440;
wire n_25441;
wire n_25442;
wire n_25443;
wire n_25444;
wire n_25445;
wire n_25446;
wire n_25447;
wire n_25448;
wire n_25449;
wire n_25450;
wire n_25451;
wire n_25452;
wire n_25453;
wire n_25454;
wire n_25455;
wire n_25456;
wire n_25457;
wire n_25458;
wire n_25459;
wire n_25460;
wire n_25461;
wire n_25462;
wire n_25463;
wire n_25464;
wire n_25465;
wire n_25466;
wire n_25467;
wire n_25468;
wire n_25469;
wire n_25470;
wire n_25471;
wire n_25472;
wire n_25473;
wire n_25474;
wire n_25475;
wire n_25476;
wire n_25477;
wire n_25478;
wire n_25479;
wire n_25480;
wire n_25481;
wire n_25482;
wire n_25483;
wire n_25484;
wire n_25485;
wire n_25486;
wire n_25487;
wire n_25488;
wire n_25489;
wire n_25490;
wire n_25491;
wire n_25492;
wire n_25493;
wire n_25494;
wire n_25495;
wire n_25496;
wire n_25497;
wire n_25498;
wire n_25499;
wire n_25500;
wire n_25501;
wire n_25502;
wire n_25503;
wire n_25504;
wire n_25505;
wire n_25506;
wire n_25507;
wire n_25508;
wire n_25509;
wire n_25510;
wire n_25511;
wire n_25512;
wire n_25513;
wire n_25514;
wire n_25515;
wire n_25516;
wire n_25517;
wire n_25518;
wire n_25519;
wire n_25520;
wire n_25521;
wire n_25522;
wire n_25523;
wire n_25524;
wire n_25525;
wire n_25526;
wire n_25527;
wire n_25528;
wire n_25529;
wire n_25530;
wire n_25531;
wire n_25532;
wire n_25533;
wire n_25534;
wire n_25535;
wire n_25536;
wire n_25537;
wire n_25538;
wire n_25539;
wire n_25540;
wire n_25541;
wire n_25542;
wire n_25543;
wire n_25544;
wire n_25545;
wire n_25546;
wire n_25547;
wire n_25548;
wire n_25549;
wire n_25550;
wire n_25551;
wire n_25552;
wire n_25553;
wire n_25554;
wire n_25555;
wire n_25556;
wire n_25557;
wire n_25558;
wire n_25559;
wire n_25560;
wire n_25561;
wire n_25562;
wire n_25563;
wire n_25564;
wire n_25565;
wire n_25566;
wire n_25567;
wire n_25568;
wire n_25569;
wire n_25570;
wire n_25571;
wire n_25572;
wire n_25573;
wire n_25574;
wire n_25575;
wire n_25576;
wire n_25577;
wire n_25578;
wire n_25579;
wire n_25580;
wire n_25581;
wire n_25582;
wire n_25583;
wire n_25584;
wire n_25585;
wire n_25586;
wire n_25587;
wire n_25588;
wire n_25589;
wire n_25590;
wire n_25591;
wire n_25592;
wire n_25593;
wire n_25594;
wire n_25595;
wire n_25596;
wire n_25597;
wire n_25598;
wire n_25599;
wire n_25600;
wire n_25601;
wire n_25602;
wire n_25603;
wire n_25604;
wire n_25605;
wire n_25606;
wire n_25607;
wire n_25608;
wire n_25609;
wire n_25610;
wire n_25611;
wire n_25612;
wire n_25613;
wire n_25614;
wire n_25615;
wire n_25616;
wire n_25617;
wire n_25618;
wire n_25619;
wire n_25620;
wire n_25621;
wire n_25622;
wire n_25623;
wire n_25624;
wire n_25625;
wire n_25626;
wire n_25627;
wire n_25628;
wire n_25629;
wire n_25630;
wire n_25631;
wire n_25632;
wire n_25633;
wire n_25634;
wire n_25635;
wire n_25636;
wire n_25637;
wire n_25638;
wire n_25639;
wire n_25640;
wire n_25641;
wire n_25642;
wire n_25643;
wire n_25644;
wire n_25645;
wire n_25646;
wire n_25647;
wire n_25648;
wire n_25649;
wire n_25650;
wire n_25651;
wire n_25652;
wire n_25653;
wire n_25654;
wire n_25655;
wire n_25656;
wire n_25657;
wire n_25658;
wire n_25659;
wire n_25660;
wire n_25661;
wire n_25662;
wire n_25663;
wire n_25664;
wire n_25665;
wire n_25666;
wire n_25667;
wire n_25668;
wire n_25669;
wire n_25670;
wire n_25671;
wire n_25672;
wire n_25673;
wire n_25674;
wire n_25675;
wire n_25676;
wire n_25677;
wire n_25678;
wire n_25679;
wire n_25680;
wire n_25681;
wire n_25682;
wire n_25683;
wire n_25684;
wire n_25685;
wire n_25686;
wire n_25687;
wire n_25688;
wire n_25689;
wire n_25690;
wire n_25691;
wire n_25692;
wire n_25693;
wire n_25694;
wire n_25695;
wire n_25696;
wire n_25697;
wire n_25698;
wire n_25699;
wire n_25700;
wire n_25701;
wire n_25702;
wire n_25703;
wire n_25704;
wire n_25705;
wire n_25706;
wire n_25707;
wire n_25708;
wire n_25709;
wire n_25710;
wire n_25711;
wire n_25712;
wire n_25713;
wire n_25714;
wire n_25715;
wire n_25716;
wire n_25717;
wire n_25718;
wire n_25719;
wire n_25720;
wire n_25721;
wire n_25722;
wire n_25723;
wire n_25724;
wire n_25725;
wire n_25726;
wire n_25727;
wire n_25728;
wire n_25729;
wire n_25730;
wire n_25731;
wire n_25732;
wire n_25733;
wire n_25734;
wire n_25735;
wire n_25736;
wire n_25737;
wire n_25738;
wire n_25739;
wire n_25740;
wire n_25741;
wire n_25742;
wire n_25743;
wire n_25744;
wire n_25745;
wire n_25746;
wire n_25747;
wire n_25748;
wire n_25749;
wire n_25750;
wire n_25751;
wire n_25752;
wire n_25753;
wire n_25754;
wire n_25755;
wire n_25756;
wire n_25757;
wire n_25758;
wire n_25759;
wire n_25760;
wire n_25761;
wire n_25762;
wire n_25763;
wire n_25764;
wire n_25765;
wire n_25766;
wire n_25767;
wire n_25768;
wire n_25769;
wire n_25770;
wire n_25771;
wire n_25772;
wire n_25773;
wire n_25774;
wire n_25775;
wire n_25776;
wire n_25777;
wire n_25778;
wire n_25779;
wire n_25780;
wire n_25781;
wire n_25782;
wire n_25783;
wire n_25784;
wire n_25785;
wire n_25786;
wire n_25787;
wire n_25788;
wire n_25789;
wire n_25790;
wire n_25791;
wire n_25792;
wire n_25793;
wire n_25794;
wire n_25795;
wire n_25796;
wire n_25797;
wire n_25798;
wire n_25799;
wire n_25800;
wire n_25801;
wire n_25802;
wire n_25803;
wire n_25804;
wire n_25805;
wire n_25806;
wire n_25807;
wire n_25808;
wire n_25809;
wire n_25810;
wire n_25811;
wire n_25812;
wire n_25813;
wire n_25814;
wire n_25815;
wire n_25816;
wire n_25817;
wire n_25818;
wire n_25819;
wire n_25820;
wire n_25821;
wire n_25822;
wire n_25823;
wire n_25824;
wire n_25825;
wire n_25826;
wire n_25827;
wire n_25828;
wire n_25829;
wire n_25830;
wire n_25831;
wire n_25832;
wire n_25833;
wire n_25834;
wire n_25835;
wire n_25836;
wire n_25837;
wire n_25838;
wire n_25839;
wire n_25840;
wire n_25841;
wire n_25842;
wire n_25843;
wire n_25844;
wire n_25845;
wire n_25846;
wire n_25847;
wire n_25848;
wire n_25849;
wire n_25850;
wire n_25851;
wire n_25852;
wire n_25853;
wire n_25854;
wire n_25855;
wire n_25856;
wire n_25857;
wire n_25858;
wire n_25859;
wire n_25860;
wire n_25861;
wire n_25862;
wire n_25863;
wire n_25864;
wire n_25865;
wire n_25866;
wire n_25867;
wire n_25868;
wire n_25869;
wire n_25870;
wire n_25871;
wire n_25872;
wire n_25873;
wire n_25874;
wire n_25875;
wire n_25876;
wire n_25877;
wire n_25878;
wire n_25879;
wire n_25880;
wire n_25881;
wire n_25882;
wire n_25883;
wire n_25884;
wire n_25885;
wire n_25886;
wire n_25887;
wire n_25888;
wire n_25889;
wire n_25890;
wire n_25891;
wire n_25892;
wire n_25893;
wire n_25894;
wire n_25895;
wire n_25896;
wire n_25897;
wire n_25898;
wire n_25899;
wire n_25900;
wire n_25901;
wire n_25902;
wire n_25903;
wire n_25904;
wire n_25905;
wire n_25906;
wire n_25907;
wire n_25908;
wire n_25909;
wire n_25910;
wire n_25911;
wire n_25912;
wire n_25913;
wire n_25914;
wire n_25915;
wire n_25916;
wire n_25917;
wire n_25918;
wire n_25919;
wire n_25920;
wire n_25921;
wire n_25922;
wire n_25923;
wire n_25924;
wire n_25925;
wire n_25926;
wire n_25927;
wire n_25928;
wire n_25929;
wire n_25930;
wire n_25931;
wire n_25932;
wire n_25933;
wire n_25934;
wire n_25935;
wire n_25936;
wire n_25937;
wire n_25938;
wire n_25939;
wire n_25940;
wire n_25941;
wire n_25942;
wire n_25943;
wire n_25944;
wire n_25945;
wire n_25946;
wire n_25947;
wire n_25948;
wire n_25949;
wire n_25950;
wire n_25951;
wire n_25952;
wire n_25953;
wire n_25954;
wire n_25955;
wire n_25956;
wire n_25957;
wire n_25958;
wire n_25959;
wire n_25960;
wire n_25961;
wire n_25962;
wire n_25963;
wire n_25964;
wire n_25965;
wire n_25966;
wire n_25967;
wire n_25968;
wire n_25969;
wire n_25970;
wire n_25971;
wire n_25972;
wire n_25973;
wire n_25974;
wire n_25975;
wire n_25976;
wire n_25977;
wire n_25978;
wire n_25979;
wire n_25980;
wire n_25981;
wire n_25982;
wire n_25983;
wire n_25984;
wire n_25985;
wire n_25986;
wire n_25987;
wire n_25988;
wire n_25989;
wire n_25990;
wire n_25991;
wire n_25992;
wire n_25993;
wire n_25994;
wire n_25995;
wire n_25996;
wire n_25997;
wire n_25998;
wire n_25999;
wire n_26000;
wire n_26001;
wire n_26002;
wire n_26003;
wire n_26004;
wire n_26005;
wire n_26006;
wire n_26007;
wire n_26008;
wire n_26009;
wire n_26010;
wire n_26011;
wire n_26012;
wire n_26013;
wire n_26014;
wire n_26015;
wire n_26016;
wire n_26017;
wire n_26018;
wire n_26019;
wire n_26020;
wire n_26021;
wire n_26022;
wire n_26023;
wire n_26024;
wire n_26025;
wire n_26026;
wire n_26027;
wire n_26028;
wire n_26029;
wire n_26030;
wire n_26031;
wire n_26032;
wire n_26033;
wire n_26034;
wire n_26035;
wire n_26036;
wire n_26037;
wire n_26038;
wire n_26039;
wire n_26040;
wire n_26041;
wire n_26042;
wire n_26043;
wire n_26044;
wire n_26045;
wire n_26046;
wire n_26047;
wire n_26048;
wire n_26049;
wire n_26050;
wire n_26051;
wire n_26052;
wire n_26053;
wire n_26054;
wire n_26055;
wire n_26056;
wire n_26057;
wire n_26058;
wire n_26059;
wire n_26060;
wire n_26061;
wire n_26062;
wire n_26063;
wire n_26064;
wire n_26065;
wire n_26066;
wire n_26067;
wire n_26068;
wire n_26069;
wire n_26070;
wire n_26071;
wire n_26072;
wire n_26073;
wire n_26074;
wire n_26075;
wire n_26076;
wire n_26077;
wire n_26078;
wire n_26079;
wire n_26080;
wire n_26081;
wire n_26082;
wire n_26083;
wire n_26084;
wire n_26085;
wire n_26086;
wire n_26087;
wire n_26088;
wire n_26089;
wire n_26090;
wire n_26091;
wire n_26092;
wire n_26093;
wire n_26094;
wire n_26095;
wire n_26096;
wire n_26097;
wire n_26098;
wire n_26099;
wire n_26100;
wire n_26101;
wire n_26102;
wire n_26103;
wire n_26104;
wire n_26105;
wire n_26106;
wire n_26107;
wire n_26108;
wire n_26109;
wire n_26110;
wire n_26111;
wire n_26112;
wire n_26113;
wire n_26114;
wire n_26115;
wire n_26116;
wire n_26117;
wire n_26118;
wire n_26119;
wire n_26120;
wire n_26121;
wire n_26122;
wire n_26123;
wire n_26124;
wire n_26125;
wire n_26126;
wire n_26127;
wire n_26128;
wire n_26129;
wire n_26130;
wire n_26131;
wire n_26132;
wire n_26133;
wire n_26134;
wire n_26135;
wire n_26136;
wire n_26137;
wire n_26138;
wire n_26139;
wire n_26140;
wire n_26141;
wire n_26142;
wire n_26143;
wire n_26144;
wire n_26145;
wire n_26146;
wire n_26147;
wire n_26148;
wire n_26149;
wire n_26150;
wire n_26151;
wire n_26152;
wire n_26153;
wire n_26154;
wire n_26155;
wire n_26156;
wire n_26157;
wire n_26158;
wire n_26159;
wire n_26160;
wire n_26161;
wire n_26162;
wire n_26163;
wire n_26164;
wire n_26165;
wire n_26166;
wire n_26167;
wire n_26168;
wire n_26169;
wire n_26170;
wire n_26171;
wire n_26172;
wire n_26173;
wire n_26174;
wire n_26175;
wire n_26176;
wire n_26177;
wire n_26178;
wire n_26179;
wire n_26180;
wire n_26181;
wire n_26182;
wire n_26183;
wire n_26184;
wire n_26185;
wire n_26186;
wire n_26187;
wire n_26188;
wire n_26189;
wire n_26190;
wire n_26191;
wire n_26192;
wire n_26193;
wire n_26194;
wire n_26195;
wire n_26196;
wire n_26197;
wire n_26198;
wire n_26199;
wire n_26200;
wire n_26201;
wire n_26202;
wire n_26203;
wire n_26204;
wire n_26205;
wire n_26206;
wire n_26207;
wire n_26208;
wire n_26209;
wire n_26210;
wire n_26211;
wire n_26212;
wire n_26213;
wire n_26214;
wire n_26215;
wire n_26216;
wire n_26217;
wire n_26218;
wire n_26219;
wire n_26220;
wire n_26221;
wire n_26222;
wire n_26223;
wire n_26224;
wire n_26225;
wire n_26226;
wire n_26227;
wire n_26228;
wire n_26229;
wire n_26230;
wire n_26231;
wire n_26232;
wire n_26233;
wire n_26234;
wire n_26235;
wire n_26236;
wire n_26237;
wire n_26238;
wire n_26239;
wire n_26240;
wire n_26241;
wire n_26242;
wire n_26243;
wire n_26244;
wire n_26245;
wire n_26246;
wire n_26247;
wire n_26248;
wire n_26249;
wire n_26250;
wire n_26251;
wire n_26252;
wire n_26253;
wire n_26254;
wire n_26255;
wire n_26256;
wire n_26257;
wire n_26258;
wire n_26259;
wire n_26260;
wire n_26261;
wire n_26262;
wire n_26263;
wire n_26264;
wire n_26265;
wire n_26266;
wire n_26267;
wire n_26268;
wire n_26269;
wire n_26270;
wire n_26271;
wire n_26272;
wire n_26273;
wire n_26274;
wire n_26275;
wire n_26276;
wire n_26277;
wire n_26278;
wire n_26279;
wire n_26280;
wire n_26281;
wire n_26282;
wire n_26283;
wire n_26284;
wire n_26285;
wire n_26286;
wire n_26287;
wire n_26288;
wire n_26289;
wire n_26290;
wire n_26291;
wire n_26292;
wire n_26293;
wire n_26294;
wire n_26295;
wire n_26296;
wire n_26297;
wire n_26298;
wire n_26299;
wire n_26300;
wire n_26301;
wire n_26302;
wire n_26303;
wire n_26304;
wire n_26305;
wire n_26306;
wire n_26307;
wire n_26308;
wire n_26309;
wire n_26310;
wire n_26311;
wire n_26312;
wire n_26313;
wire n_26314;
wire n_26315;
wire n_26316;
wire n_26317;
wire n_26318;
wire n_26319;
wire n_26320;
wire n_26321;
wire n_26322;
wire n_26323;
wire n_26324;
wire n_26325;
wire n_26326;
wire n_26327;
wire n_26328;
wire n_26329;
wire n_26330;
wire n_26331;
wire n_26332;
wire n_26333;
wire n_26334;
wire n_26335;
wire n_26336;
wire n_26337;
wire n_26338;
wire n_26339;
wire n_26340;
wire n_26341;
wire n_26342;
wire n_26343;
wire n_26344;
wire n_26345;
wire n_26346;
wire n_26347;
wire n_26348;
wire n_26349;
wire n_26350;
wire n_26351;
wire n_26352;
wire n_26353;
wire n_26354;
wire n_26355;
wire n_26356;
wire n_26357;
wire n_26358;
wire n_26359;
wire n_26360;
wire n_26361;
wire n_26362;
wire n_26363;
wire n_26364;
wire n_26365;
wire n_26366;
wire n_26367;
wire n_26368;
wire n_26369;
wire n_26370;
wire n_26371;
wire n_26372;
wire n_26373;
wire n_26374;
wire n_26375;
wire n_26376;
wire n_26377;
wire n_26378;
wire n_26379;
wire n_26380;
wire n_26381;
wire n_26382;
wire n_26383;
wire n_26384;
wire n_26385;
wire n_26386;
wire n_26387;
wire n_26388;
wire n_26389;
wire n_26390;
wire n_26391;
wire n_26392;
wire n_26393;
wire n_26394;
wire n_26395;
wire n_26396;
wire n_26397;
wire n_26398;
wire n_26399;
wire n_26400;
wire n_26401;
wire n_26402;
wire n_26403;
wire n_26404;
wire n_26405;
wire n_26406;
wire n_26407;
wire n_26408;
wire n_26409;
wire n_26410;
wire n_26411;
wire n_26412;
wire n_26413;
wire n_26414;
wire n_26415;
wire n_26416;
wire n_26417;
wire n_26418;
wire n_26419;
wire n_26420;
wire n_26421;
wire n_26422;
wire n_26423;
wire n_26424;
wire n_26425;
wire n_26426;
wire n_26427;
wire n_26428;
wire n_26429;
wire n_26430;
wire n_26431;
wire n_26432;
wire n_26433;
wire n_26434;
wire n_26435;
wire n_26436;
wire n_26437;
wire n_26438;
wire n_26439;
wire n_26440;
wire n_26441;
wire n_26442;
wire n_26443;
wire n_26444;
wire n_26445;
wire n_26446;
wire n_26447;
wire n_26448;
wire n_26449;
wire n_26450;
wire n_26451;
wire n_26452;
wire n_26453;
wire n_26454;
wire n_26455;
wire n_26456;
wire n_26457;
wire n_26458;
wire n_26459;
wire n_26460;
wire n_26461;
wire n_26462;
wire n_26463;
wire n_26464;
wire n_26465;
wire n_26466;
wire n_26467;
wire n_26468;
wire n_26469;
wire n_26470;
wire n_26471;
wire n_26472;
wire n_26473;
wire n_26474;
wire n_26475;
wire n_26476;
wire n_26477;
wire n_26478;
wire n_26479;
wire n_26480;
wire n_26481;
wire n_26482;
wire n_26483;
wire n_26484;
wire n_26485;
wire n_26486;
wire n_26487;
wire n_26488;
wire n_26489;
wire n_26490;
wire n_26491;
wire n_26492;
wire n_26493;
wire n_26494;
wire n_26495;
wire n_26496;
wire n_26497;
wire n_26498;
wire n_26499;
wire n_26500;
wire n_26501;
wire n_26502;
wire n_26503;
wire n_26504;
wire n_26505;
wire n_26506;
wire n_26507;
wire n_26508;
wire n_26509;
wire n_26510;
wire n_26511;
wire n_26512;
wire n_26513;
wire n_26514;
wire n_26515;
wire n_26516;
wire n_26517;
wire n_26518;
wire n_26519;
wire n_26520;
wire n_26521;
wire n_26522;
wire n_26523;
wire n_26524;
wire n_26525;
wire n_26526;
wire n_26527;
wire n_26528;
wire n_26529;
wire n_26530;
wire n_26531;
wire n_26532;
wire n_26533;
wire n_26534;
wire n_26535;
wire n_26536;
wire n_26537;
wire n_26538;
wire n_26539;
wire n_26540;
wire n_26541;
wire n_26542;
wire n_26543;
wire n_26544;
wire n_26545;
wire n_26546;
wire n_26547;
wire n_26548;
wire n_26549;
wire n_26550;
wire n_26551;
wire n_26552;
wire n_26553;
wire n_26554;
wire n_26555;
wire n_26556;
wire n_26557;
wire n_26558;
wire n_26559;
wire n_26560;
wire n_26561;
wire n_26562;
wire n_26563;
wire n_26564;
wire n_26565;
wire n_26566;
wire n_26567;
wire n_26568;
wire n_26569;
wire n_26570;
wire n_26571;
wire n_26572;
wire n_26573;
wire n_26574;
wire n_26575;
wire n_26576;
wire n_26577;
wire n_26578;
wire n_26579;
wire n_26580;
wire n_26581;
wire n_26582;
wire n_26583;
wire n_26584;
wire n_26585;
wire n_26586;
wire n_26587;
wire n_26588;
wire n_26589;
wire n_26590;
wire n_26591;
wire n_26592;
wire n_26593;
wire n_26594;
wire n_26595;
wire n_26596;
wire n_26597;
wire n_26598;
wire n_26599;
wire n_26600;
wire n_26601;
wire n_26602;
wire n_26603;
wire n_26604;
wire n_26605;
wire n_26606;
wire n_26607;
wire n_26608;
wire n_26609;
wire n_26610;
wire n_26611;
wire n_26612;
wire n_26613;
wire n_26614;
wire n_26615;
wire n_26616;
wire n_26617;
wire n_26618;
wire n_26619;
wire n_26620;
wire n_26621;
wire n_26622;
wire n_26623;
wire n_26624;
wire n_26625;
wire n_26626;
wire n_26627;
wire n_26628;
wire n_26629;
wire n_26630;
wire n_26631;
wire n_26632;
wire n_26633;
wire n_26634;
wire n_26635;
wire n_26636;
wire n_26637;
wire n_26638;
wire n_26639;
wire n_26640;
wire n_26641;
wire n_26642;
wire n_26643;
wire n_26644;
wire n_26645;
wire n_26646;
wire n_26647;
wire n_26648;
wire n_26649;
wire n_26650;
wire n_26651;
wire n_26652;
wire n_26653;
wire n_26654;
wire n_26655;
wire n_26656;
wire n_26657;
wire n_26658;
wire n_26659;
wire n_26660;
wire n_26661;
wire n_26662;
wire n_26663;
wire n_26664;
wire n_26665;
wire n_26666;
wire n_26667;
wire n_26668;
wire n_26669;
wire n_26670;
wire n_26671;
wire n_26672;
wire n_26673;
wire n_26674;
wire n_26675;
wire n_26676;
wire n_26677;
wire n_26678;
wire n_26679;
wire n_26680;
wire n_26681;
wire n_26682;
wire n_26683;
wire n_26684;
wire n_26685;
wire n_26686;
wire n_26687;
wire n_26688;
wire n_26689;
wire n_26690;
wire n_26691;
wire n_26692;
wire n_26693;
wire n_26694;
wire n_26695;
wire n_26696;
wire n_26697;
wire n_26698;
wire n_26699;
wire n_26700;
wire n_26701;
wire n_26702;
wire n_26703;
wire n_26704;
wire n_26705;
wire n_26706;
wire n_26707;
wire n_26708;
wire n_26709;
wire n_26710;
wire n_26711;
wire n_26712;
wire n_26713;
wire n_26714;
wire n_26715;
wire n_26716;
wire n_26717;
wire n_26718;
wire n_26719;
wire n_26720;
wire n_26721;
wire n_26722;
wire n_26723;
wire n_26724;
wire n_26725;
wire n_26726;
wire n_26727;
wire n_26728;
wire n_26729;
wire n_26730;
wire n_26731;
wire n_26732;
wire n_26733;
wire n_26734;
wire n_26735;
wire n_26736;
wire n_26737;
wire n_26738;
wire n_26739;
wire n_26740;
wire n_26741;
wire n_26742;
wire n_26743;
wire n_26744;
wire n_26745;
wire n_26746;
wire n_26747;
wire n_26748;
wire n_26749;
wire n_26750;
wire n_26751;
wire n_26752;
wire n_26753;
wire n_26754;
wire n_26755;
wire n_26756;
wire n_26757;
wire n_26758;
wire n_26759;
wire n_26760;
wire n_26761;
wire n_26762;
wire n_26763;
wire n_26764;
wire n_26765;
wire n_26766;
wire n_26767;
wire n_26768;
wire n_26769;
wire n_26770;
wire n_26771;
wire n_26772;
wire n_26773;
wire n_26774;
wire n_26775;
wire n_26776;
wire n_26777;
wire n_26778;
wire n_26779;
wire n_26780;
wire n_26781;
wire n_26782;
wire n_26783;
wire n_26784;
wire n_26785;
wire n_26786;
wire n_26787;
wire n_26788;
wire n_26789;
wire n_26790;
wire n_26791;
wire n_26792;
wire n_26793;
wire n_26794;
wire n_26795;
wire n_26796;
wire n_26797;
wire n_26798;
wire n_26799;
wire n_26800;
wire n_26801;
wire n_26802;
wire n_26803;
wire n_26804;
wire n_26805;
wire n_26806;
wire n_26807;
wire n_26808;
wire n_26809;
wire n_26810;
wire n_26811;
wire n_26812;
wire n_26813;
wire n_26814;
wire n_26815;
wire n_26816;
wire n_26817;
wire n_26818;
wire n_26819;
wire n_26820;
wire n_26821;
wire n_26822;
wire n_26823;
wire n_26824;
wire n_26825;
wire n_26826;
wire n_26827;
wire n_26828;
wire n_26829;
wire n_26830;
wire n_26831;
wire n_26832;
wire n_26833;
wire n_26834;
wire n_26835;
wire n_26836;
wire n_26837;
wire n_26838;
wire n_26839;
wire n_26840;
wire n_26841;
wire n_26842;
wire n_26843;
wire n_26844;
wire n_26845;
wire n_26846;
wire n_26847;
wire n_26848;
wire n_26849;
wire n_26850;
wire n_26851;
wire n_26852;
wire n_26853;
wire n_26854;
wire n_26855;
wire n_26856;
wire n_26857;
wire n_26858;
wire n_26859;
wire n_26860;
wire n_26861;
wire n_26862;
wire n_26863;
wire n_26864;
wire n_26865;
wire n_26866;
wire n_26867;
wire n_26868;
wire n_26869;
wire n_26870;
wire n_26871;
wire n_26872;
wire n_26873;
wire n_26874;
wire n_26875;
wire n_26876;
wire n_26877;
wire n_26878;
wire n_26879;
wire n_26880;
wire n_26881;
wire n_26882;
wire n_26883;
wire n_26884;
wire n_26885;
wire n_26886;
wire n_26887;
wire n_26888;
wire n_26889;
wire n_26890;
wire n_26891;
wire n_26892;
wire n_26893;
wire n_26894;
wire n_26895;
wire n_26896;
wire n_26897;
wire n_26898;
wire n_26899;
wire n_26900;
wire n_26901;
wire n_26902;
wire n_26903;
wire n_26904;
wire n_26905;
wire n_26906;
wire n_26907;
wire n_26908;
wire n_26909;
wire n_26910;
wire n_26911;
wire n_26912;
wire n_26913;
wire n_26914;
wire n_26915;
wire n_26916;
wire n_26917;
wire n_26918;
wire n_26919;
wire n_26920;
wire n_26921;
wire n_26922;
wire n_26923;
wire n_26924;
wire n_26925;
wire n_26926;
wire n_26927;
wire n_26928;
wire n_26929;
wire n_26930;
wire n_26931;
wire n_26932;
wire n_26933;
wire n_26934;
wire n_26935;
wire n_26936;
wire n_26937;
wire n_26938;
wire n_26939;
wire n_26940;
wire n_26941;
wire n_26942;
wire n_26943;
wire n_26944;
wire n_26945;
wire n_26946;
wire n_26947;
wire n_26948;
wire n_26949;
wire n_26950;
wire n_26951;
wire n_26952;
wire n_26953;
wire n_26954;
wire n_26955;
wire n_26956;
wire n_26957;
wire n_26958;
wire n_26959;
wire n_26960;
wire n_26961;
wire n_26962;
wire n_26963;
wire n_26964;
wire n_26965;
wire n_26966;
wire n_26967;
wire n_26968;
wire n_26969;
wire n_26970;
wire n_26971;
wire n_26972;
wire n_26973;
wire n_26974;
wire n_26975;
wire n_26976;
wire n_26977;
wire n_26978;
wire n_26979;
wire n_26980;
wire n_26981;
wire n_26982;
wire n_26983;
wire n_26984;
wire n_26985;
wire n_26986;
wire n_26987;
wire n_26988;
wire n_26989;
wire n_26990;
wire n_26991;
wire n_26992;
wire n_26993;
wire n_26994;
wire n_26995;
wire n_26996;
wire n_26997;
wire n_26998;
wire n_26999;
wire n_27000;
wire n_27001;
wire n_27002;
wire n_27003;
wire n_27004;
wire n_27005;
wire n_27006;
wire n_27007;
wire n_27008;
wire n_27009;
wire n_27010;
wire n_27011;
wire n_27012;
wire n_27013;
wire n_27014;
wire n_27015;
wire n_27016;
wire n_27017;
wire n_27018;
wire n_27019;
wire n_27020;
wire n_27021;
wire n_27022;
wire n_27023;
wire n_27024;
wire n_27025;
wire n_27026;
wire n_27027;
wire n_27028;
wire n_27029;
wire n_27030;
wire n_27031;
wire n_27032;
wire n_27033;
wire n_27034;
wire n_27035;
wire n_27036;
wire n_27037;
wire n_27038;
wire n_27039;
wire n_27040;
wire n_27041;
wire n_27042;
wire n_27043;
wire n_27044;
wire n_27045;
wire n_27046;
wire n_27047;
wire n_27048;
wire n_27049;
wire n_27050;
wire n_27051;
wire n_27052;
wire n_27053;
wire n_27054;
wire n_27055;
wire n_27056;
wire n_27057;
wire n_27058;
wire n_27059;
wire n_27060;
wire n_27061;
wire n_27062;
wire n_27063;
wire n_27064;
wire n_27065;
wire n_27066;
wire n_27067;
wire n_27068;
wire n_27069;
wire n_27070;
wire n_27071;
wire n_27072;
wire n_27073;
wire n_27074;
wire n_27075;
wire n_27076;
wire n_27077;
wire n_27078;
wire n_27079;
wire n_27080;
wire n_27081;
wire n_27082;
wire n_27083;
wire n_27084;
wire n_27085;
wire n_27086;
wire n_27087;
wire n_27088;
wire n_27089;
wire n_27090;
wire n_27091;
wire n_27092;
wire n_27093;
wire n_27094;
wire n_27095;
wire n_27096;
wire n_27097;
wire n_27098;
wire n_27099;
wire n_27100;
wire n_27101;
wire n_27102;
wire n_27103;
wire n_27104;
wire n_27105;
wire n_27106;
wire n_27107;
wire n_27108;
wire n_27109;
wire n_27110;
wire n_27111;
wire n_27112;
wire n_27113;
wire n_27114;
wire n_27115;
wire n_27116;
wire n_27117;
wire n_27118;
wire n_27119;
wire n_27120;
wire n_27121;
wire n_27122;
wire n_27123;
wire n_27124;
wire n_27125;
wire n_27126;
wire n_27127;
wire n_27128;
wire n_27129;
wire n_27130;
wire n_27131;
wire n_27132;
wire n_27133;
wire n_27134;
wire n_27135;
wire n_27136;
wire n_27137;
wire n_27138;
wire n_27139;
wire n_27140;
wire n_27141;
wire n_27142;
wire n_27143;
wire n_27144;
wire n_27145;
wire n_27146;
wire n_27147;
wire n_27148;
wire n_27149;
wire n_27150;
wire n_27151;
wire n_27152;
wire n_27153;
wire n_27154;
wire n_27155;
wire n_27156;
wire n_27157;
wire n_27158;
wire n_27159;
wire n_27160;
wire n_27161;
wire n_27162;
wire n_27163;
wire n_27164;
wire n_27165;
wire n_27166;
wire n_27167;
wire n_27168;
wire n_27169;
wire n_27170;
wire n_27171;
wire n_27172;
wire n_27173;
wire n_27174;
wire n_27175;
wire n_27176;
wire n_27177;
wire n_27178;
wire n_27179;
wire n_27180;
wire n_27181;
wire n_27182;
wire n_27183;
wire n_27184;
wire n_27185;
wire n_27186;
wire n_27187;
wire n_27188;
wire n_27189;
wire n_27190;
wire n_27191;
wire n_27192;
wire n_27193;
wire n_27194;
wire n_27195;
wire n_27196;
wire n_27197;
wire n_27198;
wire n_27199;
wire n_27200;
wire n_27201;
wire n_27202;
wire n_27203;
wire n_27204;
wire n_27205;
wire n_27206;
wire n_27207;
wire n_27208;
wire n_27209;
wire n_27210;
wire n_27211;
wire n_27212;
wire n_27213;
wire n_27214;
wire n_27215;
wire n_27216;
wire n_27217;
wire n_27218;
wire n_27219;
wire n_27220;
wire n_27221;
wire n_27222;
wire n_27223;
wire n_27224;
wire n_27225;
wire n_27226;
wire n_27227;
wire n_27228;
wire n_27229;
wire n_27230;
wire n_27231;
wire n_27232;
wire n_27233;
wire n_27234;
wire n_27235;
wire n_27236;
wire n_27237;
wire n_27238;
wire n_27239;
wire n_27240;
wire n_27241;
wire n_27242;
wire n_27243;
wire n_27244;
wire n_27245;
wire n_27246;
wire n_27247;
wire n_27248;
wire n_27249;
wire n_27250;
wire n_27251;
wire n_27252;
wire n_27253;
wire n_27254;
wire n_27255;
wire n_27256;
wire n_27257;
wire n_27258;
wire n_27259;
wire n_27260;
wire n_27261;
wire n_27262;
wire n_27263;
wire n_27264;
wire n_27265;
wire n_27266;
wire n_27267;
wire n_27268;
wire n_27269;
wire n_27270;
wire n_27271;
wire n_27272;
wire n_27273;
wire n_27274;
wire n_27275;
wire n_27276;
wire n_27277;
wire n_27278;
wire n_27279;
wire n_27280;
wire n_27281;
wire n_27282;
wire n_27283;
wire n_27284;
wire n_27285;
wire n_27286;
wire n_27287;
wire n_27288;
wire n_27289;
wire n_27290;
wire n_27291;
wire n_27292;
wire n_27293;
wire n_27294;
wire n_27295;
wire n_27296;
wire n_27297;
wire n_27298;
wire n_27299;
wire n_27300;
wire n_27301;
wire n_27302;
wire n_27303;
wire n_27304;
wire n_27305;
wire n_27306;
wire n_27307;
wire n_27308;
wire n_27309;
wire n_27310;
wire n_27311;
wire n_27312;
wire n_27313;
wire n_27314;
wire n_27315;
wire n_27316;
wire n_27317;
wire n_27318;
wire n_27319;
wire n_27320;
wire n_27321;
wire n_27322;
wire n_27323;
wire n_27324;
wire n_27325;
wire n_27326;
wire n_27327;
wire n_27328;
wire n_27329;
wire n_27330;
wire n_27331;
wire n_27332;
wire n_27333;
wire n_27334;
wire n_27335;
wire n_27336;
wire n_27337;
wire n_27338;
wire n_27339;
wire n_27340;
wire n_27341;
wire n_27342;
wire n_27343;
wire n_27344;
wire n_27345;
wire n_27346;
wire n_27347;
wire n_27348;
wire n_27349;
wire n_27350;
wire n_27351;
wire n_27352;
wire n_27353;
wire n_27354;
wire n_27355;
wire n_27356;
wire n_27357;
wire n_27358;
wire n_27359;
wire n_27360;
wire n_27361;
wire n_27362;
wire n_27363;
wire n_27364;
wire n_27365;
wire n_27366;
wire n_27367;
wire n_27368;
wire n_27369;
wire n_27370;
wire n_27371;
wire n_27372;
wire n_27373;
wire n_27374;
wire n_27375;
wire n_27376;
wire n_27377;
wire n_27378;
wire n_27379;
wire n_27380;
wire n_27381;
wire n_27382;
wire n_27383;
wire n_27384;
wire n_27385;
wire n_27386;
wire n_27387;
wire n_27388;
wire n_27389;
wire n_27390;
wire n_27391;
wire n_27392;
wire n_27393;
wire n_27394;
wire n_27395;
wire n_27396;
wire n_27397;
wire n_27398;
wire n_27399;
wire n_27400;
wire n_27401;
wire n_27402;
wire n_27403;
wire n_27404;
wire n_27405;
wire n_27406;
wire n_27407;
wire n_27408;
wire n_27409;
wire n_27410;
wire n_27411;
wire n_27412;
wire n_27413;
wire n_27414;
wire n_27415;
wire n_27416;
wire n_27417;
wire n_27418;
wire n_27419;
wire n_27420;
wire n_27421;
wire n_27422;
wire n_27423;
wire n_27424;
wire n_27425;
wire n_27426;
wire n_27427;
wire n_27428;
wire n_27429;
wire n_27430;
wire n_27431;
wire n_27432;
wire n_27433;
wire n_27434;
wire n_27435;
wire n_27436;
wire n_27437;
wire n_27438;
wire n_27439;
wire n_27440;
wire n_27441;
wire n_27442;
wire n_27443;
wire n_27444;
wire n_27445;
wire n_27446;
wire n_27447;
wire n_27448;
wire n_27449;
wire n_27450;
wire n_27451;
wire n_27452;
wire n_27453;
wire n_27454;
wire n_27455;
wire n_27456;
wire n_27457;
wire n_27458;
wire n_27459;
wire n_27460;
wire n_27461;
wire n_27462;
wire n_27463;
wire n_27464;
wire n_27465;
wire n_27466;
wire n_27467;
wire n_27468;
wire n_27469;
wire n_27470;
wire n_27471;
wire n_27472;
wire n_27473;
wire n_27474;
wire n_27475;
wire n_27476;
wire n_27477;
wire n_27478;
wire n_27479;
wire n_27480;
wire n_27481;
wire n_27482;
wire n_27483;
wire n_27484;
wire n_27485;
wire n_27486;
wire n_27487;
wire n_27488;
wire n_27489;
wire n_27490;
wire n_27491;
wire n_27492;
wire n_27493;
wire n_27494;
wire n_27495;
wire n_27496;
wire n_27497;
wire n_27498;
wire n_27499;
wire n_27500;
wire n_27501;
wire n_27502;
wire n_27503;
wire n_27504;
wire n_27505;
wire n_27506;
wire n_27507;
wire n_27508;
wire n_27509;
wire n_27510;
wire n_27511;
wire n_27512;
wire n_27513;
wire n_27514;
wire n_27515;
wire n_27516;
wire n_27517;
wire n_27518;
wire n_27519;
wire n_27520;
wire n_27521;
wire n_27522;
wire n_27523;
wire n_27524;
wire n_27525;
wire n_27526;
wire n_27527;
wire n_27528;
wire n_27529;
wire n_27530;
wire n_27531;
wire n_27532;
wire n_27533;
wire n_27534;
wire n_27535;
wire n_27536;
wire n_27537;
wire n_27538;
wire n_27539;
wire n_27540;
wire n_27541;
wire n_27542;
wire n_27543;
wire n_27544;
wire n_27545;
wire n_27546;
wire n_27547;
wire n_27548;
wire n_27549;
wire n_27550;
wire n_27551;
wire n_27552;
wire n_27553;
wire n_27554;
wire n_27555;
wire n_27556;
wire n_27557;
wire n_27558;
wire n_27559;
wire n_27560;
wire n_27561;
wire n_27562;
wire n_27563;
wire n_27564;
wire n_27565;
wire n_27566;
wire n_27567;
wire n_27568;
wire n_27569;
wire n_27570;
wire n_27571;
wire n_27572;
wire n_27573;
wire n_27574;
wire n_27575;
wire n_27576;
wire n_27577;
wire n_27578;
wire n_27579;
wire n_27580;
wire n_27581;
wire n_27582;
wire n_27583;
wire n_27584;
wire n_27585;
wire n_27586;
wire n_27587;
wire n_27588;
wire n_27589;
wire n_27590;
wire n_27591;
wire n_27592;
wire n_27593;
wire n_27594;
wire n_27595;
wire n_27596;
wire n_27597;
wire n_27598;
wire n_27599;
wire n_27600;
wire n_27601;
wire n_27602;
wire n_27603;
wire n_27604;
wire n_27605;
wire n_27606;
wire n_27607;
wire n_27608;
wire n_27609;
wire n_27610;
wire n_27611;
wire n_27612;
wire n_27613;
wire n_27614;
wire n_27615;
wire n_27616;
wire n_27617;
wire n_27618;
wire n_27619;
wire n_27620;
wire n_27621;
wire n_27622;
wire n_27623;
wire n_27624;
wire n_27625;
wire n_27626;
wire n_27627;
wire n_27628;
wire n_27629;
wire n_27630;
wire n_27631;
wire n_27632;
wire n_27633;
wire n_27634;
wire n_27635;
wire n_27636;
wire n_27637;
wire n_27638;
wire n_27639;
wire n_27640;
wire n_27641;
wire n_27642;
wire n_27643;
wire n_27644;
wire n_27645;
wire n_27646;
wire n_27647;
wire n_27648;
wire n_27649;
wire n_27650;
wire n_27651;
wire n_27652;
wire n_27653;
wire n_27654;
wire n_27655;
wire n_27656;
wire n_27657;
wire n_27658;
wire n_27659;
wire n_27660;
wire n_27661;
wire n_27662;
wire n_27663;
wire n_27664;
wire n_27665;
wire n_27666;
wire n_27667;
wire n_27668;
wire n_27669;
wire n_27670;
wire n_27671;
wire n_27672;
wire n_27673;
wire n_27674;
wire n_27675;
wire n_27676;
wire n_27677;
wire n_27678;
wire n_27679;
wire n_27680;
wire n_27681;
wire n_27682;
wire n_27683;
wire n_27684;
wire n_27685;
wire n_27686;
wire n_27687;
wire n_27688;
wire n_27689;
wire n_27690;
wire n_27691;
wire n_27692;
wire n_27693;
wire n_27694;
wire n_27695;
wire n_27696;
wire n_27697;
wire n_27698;
wire n_27699;
wire n_27700;
wire n_27701;
wire n_27702;
wire n_27703;
wire n_27704;
wire n_27705;
wire n_27706;
wire n_27707;
wire n_27708;
wire n_27709;
wire n_27710;
wire n_27711;
wire n_27712;
wire n_27713;
wire n_27714;
wire n_27715;
wire n_27716;
wire n_27717;
wire n_27718;
wire n_27719;
wire n_27720;
wire n_27721;
wire n_27722;
wire n_27723;
wire n_27724;
wire n_27725;
wire n_27726;
wire n_27727;
wire n_27728;
wire n_27729;
wire n_27730;
wire n_27731;
wire n_27732;
wire n_27733;
wire n_27734;
wire n_27735;
wire n_27736;
wire n_27737;
wire n_27738;
wire n_27739;
wire n_27740;
wire n_27741;
wire n_27742;
wire n_27743;
wire n_27744;
wire n_27745;
wire n_27746;
wire n_27747;
wire n_27748;
wire n_27749;
wire n_27750;
wire n_27751;
wire n_27752;
wire n_27753;
wire n_27754;
wire n_27755;
wire n_27756;
wire n_27757;
wire n_27758;
wire n_27759;
wire n_27760;
wire n_27761;
wire n_27762;
wire n_27763;
wire n_27764;
wire n_27765;
wire n_27766;
wire n_27767;
wire n_27768;
wire n_27769;
wire n_27770;
wire n_27771;
wire n_27772;
wire n_27773;
wire n_27774;
wire n_27775;
wire n_27776;
wire n_27777;
wire n_27778;
wire n_27779;
wire n_27780;
wire n_27781;
wire n_27782;
wire n_27783;
wire n_27784;
wire n_27785;
wire n_27786;
wire n_27787;
wire n_27788;
wire n_27789;
wire n_27790;
wire n_27791;
wire n_27792;
wire n_27793;
wire n_27794;
wire n_27795;
wire n_27796;
wire n_27797;
wire n_27798;
wire n_27799;
wire n_27800;
wire n_27801;
wire n_27802;
wire n_27803;
wire n_27804;
wire n_27805;
wire n_27806;
wire n_27807;
wire n_27808;
wire n_27809;
wire n_27810;
wire n_27811;
wire n_27812;
wire n_27813;
wire n_27814;
wire n_27815;
wire n_27816;
wire n_27817;
wire n_27818;
wire n_27819;
wire n_27820;
wire n_27821;
wire n_27822;
wire n_27823;
wire n_27824;
wire n_27825;
wire n_27826;
wire n_27827;
wire n_27828;
wire n_27829;
wire n_27830;
wire n_27831;
wire n_27832;
wire n_27833;
wire n_27834;
wire n_27835;
wire n_27836;
wire n_27837;
wire n_27838;
wire n_27839;
wire n_27840;
wire n_27841;
wire n_27842;
wire n_27843;
wire n_27844;
wire n_27845;
wire n_27846;
wire n_27847;
wire n_27848;
wire n_27849;
wire n_27850;
wire n_27851;
wire n_27852;
wire n_27853;
wire n_27854;
wire n_27855;
wire n_27856;
wire n_27857;
wire n_27858;
wire n_27859;
wire n_27860;
wire n_27861;
wire n_27862;
wire n_27863;
wire n_27864;
wire n_27865;
wire n_27866;
wire n_27867;
wire n_27868;
wire n_27869;
wire n_27870;
wire n_27871;
wire n_27872;
wire n_27873;
wire n_27874;
wire n_27875;
wire n_27876;
wire n_27877;
wire n_27878;
wire n_27879;
wire n_27880;
wire n_27881;
wire n_27882;
wire n_27883;
wire n_27884;
wire n_27885;
wire n_27886;
wire n_27887;
wire n_27888;
wire n_27889;
wire n_27890;
wire n_27891;
wire n_27892;
wire n_27893;
wire n_27894;
wire n_27895;
wire n_27896;
wire n_27897;
wire n_27898;
wire n_27899;
wire n_27900;
wire n_27901;
wire n_27902;
wire n_27903;
wire n_27904;
wire n_27905;
wire n_27906;
wire n_27907;
wire n_27908;
wire n_27909;
wire n_27910;
wire n_27911;
wire n_27912;
wire n_27913;
wire n_27914;
wire n_27915;
wire n_27916;
wire n_27917;
wire n_27918;
wire n_27919;
wire n_27920;
wire n_27921;
wire n_27922;
wire n_27923;
wire n_27924;
wire n_27925;
wire n_27926;
wire n_27927;
wire n_27928;
wire n_27929;
wire n_27930;
wire n_27931;
wire n_27932;
wire n_27933;
wire n_27934;
wire n_27935;
wire n_27936;
wire n_27937;
wire n_27938;
wire n_27939;
wire n_27940;
wire n_27941;
wire n_27942;
wire n_27943;
wire n_27944;
wire n_27945;
wire n_27946;
wire n_27947;
wire n_27948;
wire n_27949;
wire n_27950;
wire n_27951;
wire n_27952;
wire n_27953;
wire n_27954;
wire n_27955;
wire n_27956;
wire n_27957;
wire n_27958;
wire n_27959;
wire n_27960;
wire n_27961;
wire n_27962;
wire n_27963;
wire n_27964;
wire n_27965;
wire n_27966;
wire n_27967;
wire n_27968;
wire n_27969;
wire n_27970;
wire n_27971;
wire n_27972;
wire n_27973;
wire n_27974;
wire n_27975;
wire n_27976;
wire n_27977;
wire n_27978;
wire n_27979;
wire n_27980;
wire n_27981;
wire n_27982;
wire n_27983;
wire n_27984;
wire n_27985;
wire n_27986;
wire n_27987;
wire n_27988;
wire n_27989;
wire n_27990;
wire n_27991;
wire n_27992;
wire n_27993;
wire n_27994;
wire n_27995;
wire n_27996;
wire n_27997;
wire n_27998;
wire n_27999;
wire n_28000;
wire n_28001;
wire n_28002;
wire n_28003;
wire n_28004;
wire n_28005;
wire n_28006;
wire n_28007;
wire n_28008;
wire n_28009;
wire n_28010;
wire n_28011;
wire n_28012;
wire n_28013;
wire n_28014;
wire n_28015;
wire n_28016;
wire n_28017;
wire n_28018;
wire n_28019;
wire n_28020;
wire n_28021;
wire n_28022;
wire n_28023;
wire n_28024;
wire n_28025;
wire n_28026;
wire n_28027;
wire n_28028;
wire n_28029;
wire n_28030;
wire n_28031;
wire n_28032;
wire n_28033;
wire n_28034;
wire n_28035;
wire n_28036;
wire n_28037;
wire n_28038;
wire n_28039;
wire n_28040;
wire n_28041;
wire n_28042;
wire n_28043;
wire n_28044;
wire n_28045;
wire n_28046;
wire n_28047;
wire n_28048;
wire n_28049;
wire n_28050;
wire n_28051;
wire n_28052;
wire n_28053;
wire n_28054;
wire n_28055;
wire n_28056;
wire n_28057;
wire n_28058;
wire n_28059;
wire n_28060;
wire n_28061;
wire n_28062;
wire n_28063;
wire n_28064;
wire n_28065;
wire n_28066;
wire n_28067;
wire n_28068;
wire n_28069;
wire n_28070;
wire n_28071;
wire n_28072;
wire n_28073;
wire n_28074;
wire n_28075;
wire n_28076;
wire n_28077;
wire n_28078;
wire n_28079;
wire n_28080;
wire n_28081;
wire n_28082;
wire n_28083;
wire n_28084;
wire n_28085;
wire n_28086;
wire n_28087;
wire n_28088;
wire n_28089;
wire n_28090;
wire n_28091;
wire n_28092;
wire n_28093;
wire n_28094;
wire n_28095;
wire n_28096;
wire n_28097;
wire n_28098;
wire n_28099;
wire n_28100;
wire n_28101;
wire n_28102;
wire n_28103;
wire n_28104;
wire n_28105;
wire n_28106;
wire n_28107;
wire n_28108;
wire n_28109;
wire n_28110;
wire n_28111;
wire n_28112;
wire n_28113;
wire n_28114;
wire n_28115;
wire n_28116;
wire n_28117;
wire n_28118;
wire n_28119;
wire n_28120;
wire n_28121;
wire n_28122;
wire n_28123;
wire n_28124;
wire n_28125;
wire n_28126;
wire n_28127;
wire n_28128;
wire n_28129;
wire n_28130;
wire n_28131;
wire n_28132;
wire n_28133;
wire n_28134;
wire n_28135;
wire n_28136;
wire n_28137;
wire n_28138;
wire n_28139;
wire n_28140;
wire n_28141;
wire n_28142;
wire n_28143;
wire n_28144;
wire n_28145;
wire n_28146;
wire n_28147;
wire n_28148;
wire n_28149;
wire n_28150;
wire n_28151;
wire n_28152;
wire n_28153;
wire n_28154;
wire n_28155;
wire n_28156;
wire n_28157;
wire n_28158;
wire n_28159;
wire n_28160;
wire n_28161;
wire n_28162;
wire n_28163;
wire n_28164;
wire n_28165;
wire n_28166;
wire n_28167;
wire n_28168;
wire n_28169;
wire n_28170;
wire n_28171;
wire n_28172;
wire n_28173;
wire n_28174;
wire n_28175;
wire n_28176;
wire n_28177;
wire n_28178;
wire n_28179;
wire n_28180;
wire n_28181;
wire n_28182;
wire n_28183;
wire n_28184;
wire n_28185;
wire n_28186;
wire n_28187;
wire n_28188;
wire n_28189;
wire n_28190;
wire n_28191;
wire n_28192;
wire n_28193;
wire n_28194;
wire n_28195;
wire n_28196;
wire n_28197;
wire n_28198;
wire n_28199;
wire n_28200;
wire n_28201;
wire n_28202;
wire n_28203;
wire n_28204;
wire n_28205;
wire n_28206;
wire n_28207;
wire n_28208;
wire n_28209;
wire n_28210;
wire n_28211;
wire n_28212;
wire n_28213;
wire n_28214;
wire n_28215;
wire n_28216;
wire n_28217;
wire n_28218;
wire n_28219;
wire n_28220;
wire n_28221;
wire n_28222;
wire n_28223;
wire n_28224;
wire n_28225;
wire n_28226;
wire n_28227;
wire n_28228;
wire n_28229;
wire n_28230;
wire n_28231;
wire n_28232;
wire n_28233;
wire n_28234;
wire n_28235;
wire n_28236;
wire n_28237;
wire n_28238;
wire n_28239;
wire n_28240;
wire n_28241;
wire n_28242;
wire n_28243;
wire n_28244;
wire n_28245;
wire n_28246;
wire n_28247;
wire n_28248;
wire n_28249;
wire n_28250;
wire n_28251;
wire n_28252;
wire n_28253;
wire n_28254;
wire n_28255;
wire n_28256;
wire n_28257;
wire n_28258;
wire n_28259;
wire n_28260;
wire n_28261;
wire n_28262;
wire n_28263;
wire n_28264;
wire n_28265;
wire n_28266;
wire n_28267;
wire n_28268;
wire n_28269;
wire n_28270;
wire n_28271;
wire n_28272;
wire n_28273;
wire n_28274;
wire n_28275;
wire n_28276;
wire n_28277;
wire n_28278;
wire n_28279;
wire n_28280;
wire n_28281;
wire n_28282;
wire n_28283;
wire n_28284;
wire n_28285;
wire n_28286;
wire n_28287;
wire n_28288;
wire n_28289;
wire n_28290;
wire n_28291;
wire n_28292;
wire n_28293;
wire n_28294;
wire n_28295;
wire n_28296;
wire n_28297;
wire n_28298;
wire n_28299;
wire n_28300;
wire n_28301;
wire n_28302;
wire n_28303;
wire n_28304;
wire n_28305;
wire n_28306;
wire n_28307;
wire n_28308;
wire n_28309;
wire n_28310;
wire n_28311;
wire n_28312;
wire n_28313;
wire n_28314;
wire n_28315;
wire n_28316;
wire n_28317;
wire n_28318;
wire n_28319;
wire n_28320;
wire n_28321;
wire n_28322;
wire n_28323;
wire n_28324;
wire n_28325;
wire n_28326;
wire n_28327;
wire n_28328;
wire n_28329;
wire n_28330;
wire n_28331;
wire n_28332;
wire n_28333;
wire n_28334;
wire n_28335;
wire n_28336;
wire n_28337;
wire n_28338;
wire n_28339;
wire n_28340;
wire n_28341;
wire n_28342;
wire n_28343;
wire n_28344;
wire n_28345;
wire n_28346;
wire n_28347;
wire n_28348;
wire n_28349;
wire n_28350;
wire n_28351;
wire n_28352;
wire n_28353;
wire n_28354;
wire n_28355;
wire n_28356;
wire n_28357;
wire n_28358;
wire n_28359;
wire n_28360;
wire n_28361;
wire n_28362;
wire n_28363;
wire n_28364;
wire n_28365;
wire n_28366;
wire n_28367;
wire n_28368;
wire n_28369;
wire n_28370;
wire n_28371;
wire n_28372;
wire n_28373;
wire n_28374;
wire n_28375;
wire n_28376;
wire n_28377;
wire n_28378;
wire n_28379;
wire n_28380;
wire n_28381;
wire n_28382;
wire n_28383;
wire n_28384;
wire n_28385;
wire n_28386;
wire n_28387;
wire n_28388;
wire n_28389;
wire n_28390;
wire n_28391;
wire n_28392;
wire n_28393;
wire n_28394;
wire n_28395;
wire n_28396;
wire n_28397;
wire n_28398;
wire n_28399;
wire n_28400;
wire n_28401;
wire n_28402;
wire n_28403;
wire n_28404;
wire n_28405;
wire n_28406;
wire n_28407;
wire n_28408;
wire n_28409;
wire n_28410;
wire n_28411;
wire n_28412;
wire n_28413;
wire n_28414;
wire n_28415;
wire n_28416;
wire n_28417;
wire n_28418;
wire n_28419;
wire n_28420;
wire n_28421;
wire n_28422;
wire n_28423;
wire n_28424;
wire n_28425;
wire n_28426;
wire n_28427;
wire n_28428;
wire n_28429;
wire n_28430;
wire n_28431;
wire n_28432;
wire n_28433;
wire n_28434;
wire n_28435;
wire n_28436;
wire n_28437;
wire n_28438;
wire n_28439;
wire n_28440;
wire n_28441;
wire n_28442;
wire n_28443;
wire n_28444;
wire n_28445;
wire n_28446;
wire n_28447;
wire n_28448;
wire n_28449;
wire n_28450;
wire n_28451;
wire n_28452;
wire n_28453;
wire n_28454;
wire n_28455;
wire n_28456;
wire n_28457;
wire n_28458;
wire n_28459;
wire n_28460;
wire n_28461;
wire n_28462;
wire n_28463;
wire n_28464;
wire n_28465;
wire n_28466;
wire n_28467;
wire n_28468;
wire n_28469;
wire n_28470;
wire n_28471;
wire n_28472;
wire n_28473;
wire n_28474;
wire n_28475;
wire n_28476;
wire n_28477;
wire n_28478;
wire n_28479;
wire n_28480;
wire n_28481;
wire n_28482;
wire n_28483;
wire n_28484;
wire n_28485;
wire n_28486;
wire n_28487;
wire n_28488;
wire n_28489;
wire n_28490;
wire n_28491;
wire n_28492;
wire n_28493;
wire n_28494;
wire n_28495;
wire n_28496;
wire n_28497;
wire n_28498;
wire n_28499;
wire n_28500;
wire n_28501;
wire n_28502;
wire n_28503;
wire n_28504;
wire n_28505;
wire n_28506;
wire n_28507;
wire n_28508;
wire n_28509;
wire n_28510;
wire n_28511;
wire n_28512;
wire n_28513;
wire n_28514;
wire n_28515;
wire n_28516;
wire n_28517;
wire n_28518;
wire n_28519;
wire n_28520;
wire n_28521;
wire n_28522;
wire n_28523;
wire n_28524;
wire n_28525;
wire n_28526;
wire n_28527;
wire n_28528;
wire n_28529;
wire n_28530;
wire n_28531;
wire n_28532;
wire n_28533;
wire n_28534;
wire n_28535;
wire n_28536;
wire n_28537;
wire n_28538;
wire n_28539;
wire n_28540;
wire n_28541;
wire n_28542;
wire n_28543;
wire n_28544;
wire n_28545;
wire n_28546;
wire n_28547;
wire n_28548;
wire n_28549;
wire n_28550;
wire n_28551;
wire n_28552;
wire n_28553;
wire n_28554;
wire n_28555;
wire n_28556;
wire n_28557;
wire n_28558;
wire n_28559;
wire n_28560;
wire n_28561;
wire n_28562;
wire n_28563;
wire n_28564;
wire n_28565;
wire n_28566;
wire n_28567;
wire n_28568;
wire n_28569;
wire n_28570;
wire n_28571;
wire n_28572;
wire n_28573;
wire n_28574;
wire n_28575;
wire n_28576;
wire n_28577;
wire n_28578;
wire n_28579;
wire n_28580;
wire n_28581;
wire n_28582;
wire n_28583;
wire n_28584;
wire n_28585;
wire n_28586;
wire n_28587;
wire n_28588;
wire n_28589;
wire n_28590;
wire n_28591;
wire n_28592;
wire n_28593;
wire n_28594;
wire n_28595;
wire n_28596;
wire n_28597;
wire n_28598;
wire n_28599;
wire n_28600;
wire n_28601;
wire n_28602;
wire n_28603;
wire n_28604;
wire n_28605;
wire n_28606;
wire n_28607;
wire n_28608;
wire n_28609;
wire n_28610;
wire n_28611;
wire n_28612;
wire n_28613;
wire n_28614;
wire n_28615;
wire n_28616;
wire n_28617;
wire n_28618;
wire n_28619;
wire n_28620;
wire n_28621;
wire n_28622;
wire n_28623;
wire n_28624;
wire n_28625;
wire n_28626;
wire n_28627;
wire n_28628;
wire n_28629;
wire n_28630;
wire n_28631;
wire n_28632;
wire n_28633;
wire n_28634;
wire n_28635;
wire n_28636;
wire n_28637;
wire n_28638;
wire n_28639;
wire n_28640;
wire n_28641;
wire n_28642;
wire n_28643;
wire n_28644;
wire n_28645;
wire n_28646;
wire n_28647;
wire n_28648;
wire n_28649;
wire n_28650;
wire n_28651;
wire n_28652;
wire n_28653;
wire n_28654;
wire n_28655;
wire n_28656;
wire n_28657;
wire n_28658;
wire n_28659;
wire n_28660;
wire n_28661;
wire n_28662;
wire n_28663;
wire n_28664;
wire n_28665;
wire n_28666;
wire n_28667;
wire n_28668;
wire n_28669;
wire n_28670;
wire n_28671;
wire n_28672;
wire n_28673;
wire n_28674;
wire n_28675;
wire n_28676;
wire n_28677;
wire n_28678;
wire n_28679;
wire n_28680;
wire n_28681;
wire n_28682;
wire n_28683;
wire n_28684;
wire n_28685;
wire n_28686;
wire n_28687;
wire n_28688;
wire n_28689;
wire n_28690;
wire n_28691;
wire n_28692;
wire n_28693;
wire n_28694;
wire n_28695;
wire n_28696;
wire n_28697;
wire n_28698;
wire n_28699;
wire n_28700;
wire n_28701;
wire n_28702;
wire n_28703;
wire n_28704;
wire n_28705;
wire n_28706;
wire n_28707;
wire n_28708;
wire n_28709;
wire n_28710;
wire n_28711;
wire n_28712;
wire n_28713;
wire n_28714;
wire n_28715;
wire n_28716;
wire n_28717;
wire n_28718;
wire n_28719;
wire n_28720;
wire n_28721;
wire n_28722;
wire n_28723;
wire n_28724;
wire n_28725;
wire n_28726;
wire n_28727;
wire n_28728;
wire n_28729;
wire n_28730;
wire n_28731;
wire n_28732;
wire n_28733;
wire n_28734;
wire n_28735;
wire n_28736;
wire n_28737;
wire n_28738;
wire n_28739;
wire n_28740;
wire n_28741;
wire n_28742;
wire n_28743;
wire n_28744;
wire n_28745;
wire n_28746;
wire n_28747;
wire n_28748;
wire n_28749;
wire n_28750;
wire n_28751;
wire n_28752;
wire n_28753;
wire n_28754;
wire n_28755;
wire n_28756;
wire n_28757;
wire n_28758;
wire n_28759;
wire n_28760;
wire n_28761;
wire n_28762;
wire n_28763;
wire n_28764;
wire n_28765;
wire n_28766;
wire n_28767;
wire n_28768;
wire n_28769;
wire n_28770;
wire n_28771;
wire n_28772;
wire n_28773;
wire n_28774;
wire n_28775;
wire n_28776;
wire n_28777;
wire n_28778;
wire n_28779;
wire n_28780;
wire n_28781;
wire n_28782;
wire n_28783;
wire n_28784;
wire n_28785;
wire n_28786;
wire n_28787;
wire n_28788;
wire n_28789;
wire n_28790;
wire n_28791;
wire n_28792;
wire n_28793;
wire n_28794;
wire n_28795;
wire n_28796;
wire n_28797;
wire n_28798;
wire n_28799;
wire n_28800;
wire n_28801;
wire n_28802;
wire n_28803;
wire n_28804;
wire n_28805;
wire n_28806;
wire n_28807;
wire n_28808;
wire n_28809;
wire n_28810;
wire n_28811;
wire n_28812;
wire n_28813;
wire n_28814;
wire n_28815;
wire n_28816;
wire n_28817;
wire n_28818;
wire n_28819;
wire n_28820;
wire n_28821;
wire n_28822;
wire n_28823;
wire n_28824;
wire n_28825;
wire n_28826;
wire n_28827;
wire n_28828;
wire n_28829;
wire n_28830;
wire n_28831;
wire n_28832;
wire n_28833;
wire n_28834;
wire n_28835;
wire n_28836;
wire n_28837;
wire n_28838;
wire n_28839;
wire n_28840;
wire n_28841;
wire n_28842;
wire n_28843;
wire n_28844;
wire n_28845;
wire n_28846;
wire n_28847;
wire n_28848;
wire n_28849;
wire n_28850;
wire n_28851;
wire n_28852;
wire n_28853;
wire n_28854;
wire n_28855;
wire n_28856;
wire n_28857;
wire n_28858;
wire n_28859;
wire n_28860;
wire n_28861;
wire n_28862;
wire n_28863;
wire n_28864;
wire n_28865;
wire n_28866;
wire n_28867;
wire n_28868;
wire n_28869;
wire n_28870;
wire n_28871;
wire n_28872;
wire n_28873;
wire n_28874;
wire n_28875;
wire n_28876;
wire n_28877;
wire n_28878;
wire n_28879;
wire n_28880;
wire n_28881;
wire n_28882;
wire n_28883;
wire n_28884;
wire n_28885;
wire n_28886;
wire n_28887;
wire n_28888;
wire n_28889;
wire n_28890;
wire n_28891;
wire n_28892;
wire n_28893;
wire n_28894;
wire n_28895;
wire n_28896;
wire n_28897;
wire n_28898;
wire n_28899;
wire n_28900;
wire n_28901;
wire n_28902;
wire n_28903;
wire n_28904;
wire n_28905;
wire n_28906;
wire n_28907;
wire n_28908;
wire n_28909;
wire n_28910;
wire n_28911;
wire n_28912;
wire n_28913;
wire n_28914;
wire n_28915;
wire n_28916;
wire n_28917;
wire n_28918;
wire n_28919;
wire n_28920;
wire n_28921;
wire n_28922;
wire n_28923;
wire n_28924;
wire n_28925;
wire n_28926;
wire n_28927;
wire n_28928;
wire n_28929;
wire n_28930;
wire n_28931;
wire n_28932;
wire n_28933;
wire n_28934;
wire n_28935;
wire n_28936;
wire n_28937;
wire n_28938;
wire n_28939;
wire n_28940;
wire n_28941;
wire n_28942;
wire n_28943;
wire n_28944;
wire n_28945;
wire n_28946;
wire n_28947;
wire n_28948;
wire n_28949;
wire n_28950;
wire n_28951;
wire n_28952;
wire n_28953;
wire n_28954;
wire n_28955;
wire n_28956;
wire n_28957;
wire n_28958;
wire n_28959;
wire n_28960;
wire n_28961;
wire n_28962;
wire n_28963;
wire n_28964;
wire n_28965;
wire n_28966;
wire n_28967;
wire n_28968;
wire n_28969;
wire n_28970;
wire n_28971;
wire n_28972;
wire n_28973;
wire n_28974;
wire n_28975;
wire n_28976;
wire n_28977;
wire n_28978;
wire n_28979;
wire n_28980;
wire n_28981;
wire n_28982;
wire n_28983;
wire n_28984;
wire n_28985;
wire n_28986;
wire n_28987;
wire n_28988;
wire n_28989;
wire n_28990;
wire n_28991;
wire n_28992;
wire n_28993;
wire n_28994;
wire n_28995;
wire n_28996;
wire n_28997;
wire n_28998;
wire n_28999;
wire n_29000;
wire n_29001;
wire n_29002;
wire n_29003;
wire n_29004;
wire n_29005;
wire n_29006;
wire n_29007;
wire n_29008;
wire n_29009;
wire n_29010;
wire n_29011;
wire n_29012;
wire n_29013;
wire n_29014;
wire n_29015;
wire n_29016;
wire n_29017;
wire n_29018;
wire n_29019;
wire n_29020;
wire n_29021;
wire n_29022;
wire n_29023;
wire n_29024;
wire n_29025;
wire n_29026;
wire n_29027;
wire n_29028;
wire n_29029;
wire n_29030;
wire n_29031;
wire n_29032;
wire n_29033;
wire n_29034;
wire n_29035;
wire n_29036;
wire n_29037;
wire n_29038;
wire n_29039;
wire n_29040;
wire n_29041;
wire n_29042;
wire n_29043;
wire n_29044;
wire n_29045;
wire n_29046;
wire n_29047;
wire n_29048;
wire n_29049;
wire n_29050;
wire n_29051;
wire n_29052;
wire n_29053;
wire n_29054;
wire n_29055;
wire n_29056;
wire n_29057;
wire n_29058;
wire n_29059;
wire n_29060;
wire n_29061;
wire n_29062;
wire n_29063;
wire n_29064;
wire n_29065;
wire n_29066;
wire n_29067;
wire n_29068;
wire n_29069;
wire n_29070;
wire n_29071;
wire n_29072;
wire n_29073;
wire n_29074;
wire n_29075;
wire n_29076;
wire n_29077;
wire n_29078;
wire n_29079;
wire n_29080;
wire n_29081;
wire n_29082;
wire n_29083;
wire n_29084;
wire n_29085;
wire n_29086;
wire n_29087;
wire n_29088;
wire n_29089;
wire n_29090;
wire n_29091;
wire n_29092;
wire n_29093;
wire n_29094;
wire n_29095;
wire n_29096;
wire n_29097;
wire n_29098;
wire n_29099;
wire n_29100;
wire n_29101;
wire n_29102;
wire n_29103;
wire n_29104;
wire n_29105;
wire n_29106;
wire n_29107;
wire n_29108;
wire n_29109;
wire n_29110;
wire n_29111;
wire n_29112;
wire n_29113;
wire n_29114;
wire n_29115;
wire n_29116;
wire n_29117;
wire n_29118;
wire n_29119;
wire n_29120;
wire n_29121;
wire n_29122;
wire n_29123;
wire n_29124;
wire n_29125;
wire n_29126;
wire n_29127;
wire n_29128;
wire n_29129;
wire n_29130;
wire n_29131;
wire n_29132;
wire n_29133;
wire n_29134;
wire n_29135;
wire n_29136;
wire n_29137;
wire n_29138;
wire n_29139;
wire n_29140;
wire n_29141;
wire n_29142;
wire n_29143;
wire n_29144;
wire n_29145;
wire n_29146;
wire n_29147;
wire n_29148;
wire n_29149;
wire n_29150;
wire n_29151;
wire n_29152;
wire n_29153;
wire n_29154;
wire n_29155;
wire n_29156;
wire n_29157;
wire n_29158;
wire n_29159;
wire n_29160;
wire n_29161;
wire n_29162;
wire n_29163;
wire n_29164;
wire n_29165;
wire n_29166;
wire n_29167;
wire n_29168;
wire n_29169;
wire n_29170;
wire n_29171;
wire n_29172;
wire n_29173;
wire n_29174;
wire n_29175;
wire n_29176;
wire n_29177;
wire n_29178;
wire n_29179;
wire n_29180;
wire n_29181;
wire n_29182;
wire n_29183;
wire n_29184;
wire n_29185;
wire n_29186;
wire n_29187;
wire n_29188;
wire n_29189;
wire n_29190;
wire n_29191;
wire n_29192;
wire n_29193;
wire n_29194;
wire n_29195;
wire n_29196;
wire n_29197;
wire n_29198;
wire n_29199;
wire n_29200;
wire n_29201;
wire n_29202;
wire n_29203;
wire n_29204;
wire n_29205;
wire n_29206;
wire n_29207;
wire n_29208;
wire n_29209;
wire n_29210;
wire n_29211;
wire n_29212;
wire n_29213;
wire n_29214;
wire n_29215;
wire n_29216;
wire n_29217;
wire n_29218;
wire n_29219;
wire n_29220;
wire n_29221;
wire n_29222;
wire n_29223;
wire n_29224;
wire n_29225;
wire n_29226;
wire n_29227;
wire n_29228;
wire n_29229;
wire n_29230;
wire n_29231;
wire n_29232;
wire n_29233;
wire n_29234;
wire n_29235;
wire n_29236;
wire n_29237;
wire n_29238;
wire n_29239;
wire n_29240;
wire n_29241;
wire n_29242;
wire n_29243;
wire n_29244;
wire n_29245;
wire n_29246;
wire n_29247;
wire n_29248;
wire n_29249;
wire n_29250;
wire n_29251;
wire n_29252;
wire n_29253;
wire n_29254;
wire n_29255;
wire n_29256;
wire n_29257;
wire n_29258;
wire n_29259;
wire n_29260;
wire n_29261;
wire n_29262;
wire n_29263;
wire n_29264;
wire n_29265;
wire n_29266;
wire n_29267;
wire n_29268;
wire n_29269;
wire n_29270;
wire n_29271;
wire n_29272;
wire n_29273;
wire n_29274;
wire n_29275;
wire n_29276;
wire n_29277;
wire n_29278;
wire n_29279;
wire n_29280;
wire n_29281;
wire n_29282;
wire n_29283;
wire n_29284;
wire n_29285;
wire n_29286;
wire n_29287;
wire n_29288;
wire n_29289;
wire n_29290;
wire n_29291;
wire n_29292;
wire n_29293;
wire n_29294;
wire n_29295;
wire n_29296;
wire n_29297;
wire n_29298;
wire n_29299;
wire n_29300;
wire n_29301;
wire n_29302;
wire n_29303;
wire n_29304;
wire n_29305;
wire n_29306;
wire n_29307;
wire n_29308;
wire n_29309;
wire n_29310;
wire n_29311;
wire n_29312;
wire n_29313;
wire n_29314;
wire n_29315;
wire n_29316;
wire n_29317;
wire n_29318;
wire n_29319;
wire n_29320;
wire n_29321;
wire n_29322;
wire n_29323;
wire n_29324;
wire n_29325;
wire n_29326;
wire n_29327;
wire n_29328;
wire n_29329;
wire n_29330;
wire n_29331;
wire n_29332;
wire n_29333;
wire n_29334;
wire n_29335;
wire n_29336;
wire n_29337;
wire n_29338;
wire n_29339;
wire n_29340;
wire n_29341;
wire n_29342;
wire n_29343;
wire n_29344;
wire n_29345;
wire n_29346;
wire n_29347;
wire n_29348;
wire n_29349;
wire n_29350;
wire n_29351;
wire n_29352;
wire n_29353;
wire n_29354;
wire n_29355;
wire n_29356;
wire n_29357;
wire n_29358;
wire n_29359;
wire n_29360;
wire n_29361;
wire n_29362;
wire n_29363;
wire n_29364;
wire n_29365;
wire n_29366;
wire n_29367;
wire n_29368;
wire n_29369;
wire n_29370;
wire n_29371;
wire n_29372;
wire n_29373;
wire n_29374;
wire n_29375;
wire n_29376;
wire n_29377;
wire n_29378;
wire n_29379;
wire n_29380;
wire n_29381;
wire n_29382;
wire n_29383;
wire n_29384;
wire n_29385;
wire n_29386;
wire n_29387;
wire n_29388;
wire n_29389;
wire n_29390;
wire n_29391;
wire n_29392;
wire n_29393;
wire n_29394;
wire n_29395;
wire n_29396;
wire n_29397;
wire n_29398;
wire n_29399;
wire n_29400;
wire n_29401;
wire n_29402;
wire n_29403;
wire n_29404;
wire n_29405;
wire n_29406;
wire n_29407;
wire n_29408;
wire n_29409;
wire n_29410;
wire n_29411;
wire n_29412;
wire n_29413;
wire n_29414;
wire n_29415;
wire n_29416;
wire n_29417;
wire n_29418;
wire n_29419;
wire n_29420;
wire n_29421;
wire n_29422;
wire n_29423;
wire n_29424;
wire n_29425;
wire n_29426;
wire n_29427;
wire n_29428;
wire n_29429;
wire n_29430;
wire n_29431;
wire n_29432;
wire n_29433;
wire n_29434;
wire n_29435;
wire n_29436;
wire n_29437;
wire n_29438;
wire n_29439;
wire n_29440;
wire n_29441;
wire n_29442;
wire n_29443;
wire n_29444;
wire n_29445;
wire n_29446;
wire n_29447;
wire n_29448;
wire n_29449;
wire n_29450;
wire n_29451;
wire n_29452;
wire n_29453;
wire n_29454;
wire n_29455;
wire n_29456;
wire n_29457;
wire n_29458;
wire n_29459;
wire n_29460;
wire n_29461;
wire n_29462;
wire n_29463;
wire n_29464;
wire n_29465;
wire n_29466;
wire n_29467;
wire n_29468;
wire n_29469;
wire n_29470;
wire n_29471;
wire n_29472;
wire n_29473;
wire n_29474;
wire n_29475;
wire n_29476;
wire n_29477;
wire n_29478;
wire n_29479;
wire n_29480;
wire n_29481;
wire n_29482;
wire n_29483;
wire n_29484;
wire n_29485;
wire n_29486;
wire n_29487;
wire n_29488;
wire n_29489;
wire n_29490;
wire n_29491;
wire n_29492;
wire n_29493;
wire n_29494;
wire n_29495;
wire n_29496;
wire n_29497;
wire n_29498;
wire n_29499;
wire n_29500;
wire n_29501;
wire n_29502;
wire n_29503;
wire n_29504;
wire n_29505;
wire n_29506;
wire n_29507;
wire n_29508;
wire n_29509;
wire n_29510;
wire n_29511;
wire n_29512;
wire n_29513;
wire n_29514;
wire n_29515;
wire n_29516;
wire n_29517;
wire n_29518;
wire n_29519;
wire n_29520;
wire n_29521;
wire n_29522;
wire n_29523;
wire n_29524;
wire n_29525;
wire n_29526;
wire n_29527;
wire n_29528;
wire n_29529;
wire n_29530;
wire n_29531;
wire n_29532;
wire n_29533;
wire n_29534;
wire n_29535;
wire n_29536;
wire n_29537;
wire n_29538;
wire n_29539;
wire n_29540;
wire n_29541;
wire n_29542;
wire n_29543;
wire n_29544;
wire n_29545;
wire n_29546;
wire n_29547;
wire n_29548;
wire n_29549;
wire n_29550;
wire n_29551;
wire n_29552;
wire n_29553;
wire n_29554;
wire n_29555;
wire n_29556;
wire n_29557;
wire n_29558;
wire n_29559;
wire n_29560;
wire n_29561;
wire n_29562;
wire n_29563;
wire n_29564;
wire n_29565;
wire n_29566;
wire n_29567;
wire n_29568;
wire n_29569;
wire n_29570;
wire n_29571;
wire n_29572;
wire n_29573;
wire n_29574;
wire n_29575;
wire n_29576;
wire n_29577;
wire n_29578;
wire n_29579;
wire n_29580;
wire n_29581;
wire n_29582;
wire n_29583;
wire n_29584;
wire n_29585;
wire n_29586;
wire n_29587;
wire n_29588;
wire n_29589;
wire n_29590;
wire n_29591;
wire n_29592;
wire n_29593;
wire n_29594;
wire n_29595;
wire n_29596;
wire n_29597;
wire n_29598;
wire n_29599;
wire n_29600;
wire n_29601;
wire n_29602;
wire n_29603;
wire n_29604;
wire n_29605;
wire n_29606;
wire n_29607;
wire n_29608;
wire n_29609;
wire n_29610;
wire n_29611;
wire n_29612;
wire n_29613;
wire n_29614;
wire n_29615;
wire n_29616;
wire n_29617;
wire n_29618;
wire n_29619;
wire n_29620;
wire n_29621;
wire n_29622;
wire n_29623;
wire n_29624;
wire n_29625;
wire n_29626;
wire n_29627;
wire n_29628;
wire n_29629;
wire n_29630;
wire n_29631;
wire n_29632;
wire n_29633;
wire n_29634;
wire n_29635;
wire n_29636;
wire n_29637;
wire n_29638;
wire n_29639;
wire n_29640;
wire n_29641;
wire n_29642;
wire n_29643;
wire n_29644;
wire n_29645;
wire n_29646;
wire n_29647;
wire n_29648;
wire n_29649;
wire n_29650;
wire n_29651;
wire n_29652;
wire n_29653;
wire n_29654;
wire n_29655;
wire n_29656;
wire n_29657;
wire n_29658;
wire n_29659;
wire n_29660;
wire n_29661;
wire n_29662;
wire n_29663;
wire n_29664;
wire n_29665;
wire n_29666;
wire n_29667;
wire n_29668;
wire n_29669;
wire n_29670;
wire n_29671;
wire n_29672;
wire n_29673;
wire n_29674;
wire n_29675;
wire n_29676;
wire n_29677;
wire n_29678;
wire n_29679;
wire n_29680;
wire n_29681;
wire n_29682;
wire n_29683;
wire n_29684;
wire n_29685;
wire n_29686;
wire n_29687;
wire n_29688;
wire n_29689;
wire n_29690;
wire n_29691;
wire n_29692;
wire n_29693;
wire n_29694;
wire n_29695;
wire n_29696;
wire n_29697;
wire n_29698;
wire n_29699;
wire n_29700;
wire n_29701;
wire n_29702;
wire n_29703;
wire n_29704;
wire n_29705;
wire n_29706;
wire n_29707;
wire n_29708;
wire n_29709;
wire n_29710;
wire n_29711;
wire n_29712;
wire n_29713;
wire n_29714;
wire n_29715;
wire n_29716;
wire n_29717;
wire n_29718;
wire n_29719;
wire n_29720;
wire n_29721;
wire n_29722;
wire n_29723;
wire n_29724;
wire n_29725;
wire n_29726;
wire n_29727;
wire n_29728;
wire n_29729;
wire n_29730;
wire n_29731;
wire n_29732;
wire n_29733;
wire n_29734;
wire n_29735;
wire n_29736;
wire n_29737;
wire n_29738;
wire n_29739;
wire n_29740;
wire n_29741;
wire n_29742;
wire n_29743;
wire n_29744;
wire n_29745;
wire n_29746;
wire n_29747;
wire n_29748;
wire n_29749;
wire n_29750;
wire n_29751;
wire n_29752;
wire n_29753;
wire n_29754;
wire n_29755;
wire n_29756;
wire n_29757;
wire n_29758;
wire n_29759;
wire n_29760;
wire n_29761;
wire n_29762;
wire n_29763;
wire n_29764;
wire n_29765;
wire n_29766;
wire n_29767;
wire n_29768;
wire n_29769;
wire n_29770;
wire n_29771;
wire n_29772;
wire n_29773;
wire n_29774;
wire n_29775;
wire n_29776;
wire n_29777;
wire n_29778;
wire n_29779;
wire n_29780;
wire n_29781;
wire n_29782;
wire n_29783;
wire n_29784;
wire n_29785;
wire n_29786;
wire n_29787;
wire n_29788;
wire n_29789;
wire n_29790;
wire n_29791;
wire n_29792;
wire n_29793;
wire n_29794;
wire n_29795;
wire n_29796;
wire n_29797;
wire n_29798;
wire n_29799;
wire n_29800;
wire n_29801;
wire n_29802;
wire n_29803;
wire n_29804;
wire n_29805;
wire n_29806;
wire n_29807;
wire n_29808;
wire n_29809;
wire n_29810;
wire n_29811;
wire n_29812;
wire n_29813;
wire n_29814;
wire n_29815;
wire n_29816;
wire n_29817;
wire n_29818;
wire n_29819;
wire n_29820;
wire n_29821;
wire n_29822;
wire n_29823;
wire n_29824;
wire n_29825;
wire n_29826;
wire n_29827;
wire n_29828;
wire n_29829;
wire n_29830;
wire n_29831;
wire n_29832;
wire n_29833;
wire n_29834;
wire n_29835;
wire n_29836;
wire n_29837;
wire n_29838;
wire n_29839;
wire n_29840;
wire n_29841;
wire n_29842;
wire n_29843;
wire n_29844;
wire n_29845;
wire n_29846;
wire n_29847;
wire n_29848;
wire n_29849;
wire n_29850;
wire n_29851;
wire n_29852;
wire n_29853;
wire n_29854;
wire n_29855;
wire n_29856;
wire n_29857;
wire n_29858;
wire n_29859;
wire n_29860;
wire n_29861;
wire n_29862;
wire n_29863;
wire n_29864;
wire n_29865;
wire n_29866;
wire n_29867;
wire n_29868;
wire n_29869;
wire n_29870;
wire n_29871;
wire n_29872;
wire n_29873;
wire n_29874;
wire n_29875;
wire n_29876;
wire n_29877;
wire n_29878;
wire n_29879;
wire n_29880;
wire n_29881;
wire n_29882;
wire n_29883;
wire n_29884;
wire n_29885;
wire n_29886;
wire n_29887;
wire n_29888;
wire n_29889;
wire n_29890;
wire n_29891;
wire n_29892;
wire n_29893;
wire n_29894;
wire n_29895;
wire n_29896;
wire n_29897;
wire n_29898;
wire n_29899;
wire n_29900;
wire n_29901;
wire n_29902;
wire n_29903;
wire n_29904;
wire n_29905;
wire n_29906;
wire n_29907;
wire n_29908;
wire n_29909;
wire n_29910;
wire n_29911;
wire n_29912;
wire n_29913;
wire n_29914;
wire n_29915;
wire n_29916;
wire n_29917;
wire n_29918;
wire n_29919;
wire n_29920;
wire n_29921;
wire n_29922;
wire n_29923;
wire n_29924;
wire n_29925;
wire n_29926;
wire n_29927;
wire n_29928;
wire n_29929;
wire n_29930;
wire n_29931;
wire n_29932;
wire n_29933;
wire n_29934;
wire n_29935;
wire n_29936;
wire n_29937;
wire n_29938;
wire n_29939;
wire n_29940;
wire n_29941;
wire n_29942;
wire n_29943;
wire n_29944;
wire n_29945;
wire n_29946;
wire n_29947;
wire n_29948;
wire n_29949;
wire n_29950;
wire n_29951;
wire n_29952;
wire n_29953;
wire n_29954;
wire n_29955;
wire n_29956;
wire n_29957;
wire n_29958;
wire n_29959;
wire n_29960;
wire n_29961;
wire n_29962;
wire n_29963;
wire n_29964;
wire n_29965;
wire n_29966;
wire n_29967;
wire n_29968;
wire n_29969;
wire n_29970;
wire n_29971;
wire n_29972;
wire n_29973;
wire n_29974;
wire n_29975;
wire n_29976;
wire n_29977;
wire n_29978;
wire n_29979;
wire n_29980;
wire n_29981;
wire n_29982;
wire n_29983;
wire n_29984;
wire n_29985;
wire n_29986;
wire n_29987;
wire n_29988;
wire n_29989;
wire n_29990;
wire n_29991;
wire n_29992;
wire n_29993;
wire n_29994;
wire n_29995;
wire n_29996;
wire n_29997;
wire n_29998;
wire n_29999;
wire n_30000;
wire n_30001;
wire n_30002;
wire n_30003;
wire n_30004;
wire n_30005;
wire n_30006;
wire n_30007;
wire n_30008;
wire n_30009;
wire n_30010;
wire n_30011;
wire n_30012;
wire n_30013;
wire n_30014;
wire n_30015;
wire n_30016;
wire n_30017;
wire n_30018;
wire n_30019;
wire n_30020;
wire n_30021;
wire n_30022;
wire n_30023;
wire n_30024;
wire n_30025;
wire n_30026;
wire n_30027;
wire n_30028;
wire n_30029;
wire n_30030;
wire n_30031;
wire n_30032;
wire n_30033;
wire n_30034;
wire n_30035;
wire n_30036;
wire n_30037;
wire n_30038;
wire n_30039;
wire n_30040;
wire n_30041;
wire n_30042;
wire n_30043;
wire n_30044;
wire n_30045;
wire n_30046;
wire n_30047;
wire n_30048;
wire n_30049;
wire n_30050;
wire n_30051;
wire n_30052;
wire n_30053;
wire n_30054;
wire n_30055;
wire n_30056;
wire n_30057;
wire n_30058;
wire n_30059;
wire n_30060;
wire n_30061;
wire n_30062;
wire n_30063;
wire n_30064;
wire n_30065;
wire n_30066;
wire n_30067;
wire n_30068;
wire n_30069;
wire n_30070;
wire n_30071;
wire n_30072;
wire n_30073;
wire n_30074;
wire n_30075;
wire n_30076;
wire n_30077;
wire n_30078;
wire n_30079;
wire n_30080;
wire n_30081;
wire n_30082;
wire n_30083;
wire n_30084;
wire n_30085;
wire n_30086;
wire n_30087;
wire n_30088;
wire n_30089;
wire n_30090;
wire n_30091;
wire n_30092;
wire n_30093;
wire n_30094;
wire n_30095;
wire n_30096;
wire n_30097;
wire n_30098;
wire n_30099;
wire n_30100;
wire n_30101;
wire n_30102;
wire n_30103;
wire n_30104;
wire n_30105;
wire n_30106;
wire n_30107;
wire n_30108;
wire n_30109;
wire n_30110;
wire n_30111;
wire n_30112;
wire n_30113;
wire n_30114;
wire n_30115;
wire n_30116;
wire n_30117;
wire n_30118;
wire n_30119;
wire n_30120;
wire n_30121;
wire n_30122;
wire n_30123;
wire n_30124;
wire n_30125;
wire n_30126;
wire n_30127;
wire n_30128;
wire n_30129;
wire n_30130;
wire n_30131;
wire n_30132;
wire n_30133;
wire n_30134;
wire n_30135;
wire n_30136;
wire n_30137;
wire n_30138;
wire n_30139;
wire n_30140;
wire n_30141;
wire n_30142;
wire n_30143;
wire n_30144;
wire n_30145;
wire n_30146;
wire n_30147;
wire n_30148;
wire n_30149;
wire n_30150;
wire n_30151;
wire n_30152;
wire n_30153;
wire n_30154;
wire n_30155;
wire n_30156;
wire n_30157;
wire n_30158;
wire n_30159;
wire n_30160;
wire n_30161;
wire n_30162;
wire n_30163;
wire n_30164;
wire n_30165;
wire n_30166;
wire n_30167;
wire n_30168;
wire n_30169;
wire n_30170;
wire n_30171;
wire n_30172;
wire n_30173;
wire n_30174;
wire n_30175;
wire n_30176;
wire n_30177;
wire n_30178;
wire n_30179;
wire n_30180;
wire n_30181;
wire n_30182;
wire n_30183;
wire n_30184;
wire n_30185;
wire n_30186;
wire n_30187;
wire n_30188;
wire n_30189;
wire n_30190;
wire n_30191;
wire n_30192;
wire n_30193;
wire n_30194;
wire n_30195;
wire n_30196;
wire n_30197;
wire n_30198;
wire n_30199;
wire n_30200;
wire n_30201;
wire n_30202;
wire n_30203;
wire n_30204;
wire n_30205;
wire n_30206;
wire n_30207;
wire n_30208;
wire n_30209;
wire n_30210;
wire n_30211;
wire n_30212;
wire n_30213;
wire n_30214;
wire n_30215;
wire n_30216;
wire n_30217;
wire n_30218;
wire n_30219;
wire n_30220;
wire n_30221;
wire n_30222;
wire n_30223;
wire n_30224;
wire n_30225;
wire n_30226;
wire n_30227;
wire n_30228;
wire n_30229;
wire n_30230;
wire n_30231;
wire n_30232;
wire n_30233;
wire n_30234;
wire n_30235;
wire n_30236;
wire n_30237;
wire n_30238;
wire n_30239;
wire n_30240;
wire n_30241;
wire n_30242;
wire n_30243;
wire n_30244;
wire n_30245;
wire n_30246;
wire n_30247;
wire n_30248;
wire n_30249;
wire n_30250;
wire n_30251;
wire n_30252;
wire n_30253;
wire n_30254;
wire n_30255;
wire n_30256;
wire n_30257;
wire n_30258;
wire n_30259;
wire n_30260;
wire n_30261;
wire n_30262;
wire n_30263;
wire n_30264;
wire n_30265;
wire n_30266;
wire n_30267;
wire n_30268;
wire n_30269;
wire n_30270;
wire n_30271;
wire n_30272;
wire n_30273;
wire n_30274;
wire n_30275;
wire n_30276;
wire n_30277;
wire n_30278;
wire n_30279;
wire n_30280;
wire n_30281;
wire n_30282;
wire n_30283;
wire n_30284;
wire n_30285;
wire n_30286;
wire n_30287;
wire n_30288;
wire n_30289;
wire n_30290;
wire n_30291;
wire n_30292;
wire n_30293;
wire n_30294;
wire n_30295;
wire n_30296;
wire n_30297;
wire n_30298;
wire n_30299;
wire n_30300;
wire n_30301;
wire n_30302;
wire n_30303;
wire n_30304;
wire n_30305;
wire n_30306;
wire n_30307;
wire n_30308;
wire n_30309;
wire n_30310;
wire n_30311;
wire n_30312;
wire n_30313;
wire n_30314;
wire n_30315;
wire n_30316;
wire n_30317;
wire n_30318;
wire n_30319;
wire n_30320;
wire n_30321;
wire n_30322;
wire n_30323;
wire n_30324;
wire n_30325;
wire n_30326;
wire n_30327;
wire n_30328;
wire n_30329;
wire n_30330;
wire n_30331;
wire n_30332;
wire n_30333;
wire n_30334;
wire n_30335;
wire n_30336;
wire n_30337;
wire n_30338;
wire n_30339;
wire n_30340;
wire n_30341;
wire n_30342;
wire n_30343;
wire n_30344;
wire n_30345;
wire n_30346;
wire n_30347;
wire n_30348;
wire n_30349;
wire n_30350;
wire n_30351;
wire n_30352;
wire n_30353;
wire n_30354;
wire n_30355;
wire n_30356;
wire n_30357;
wire n_30358;
wire n_30359;
wire n_30360;
wire n_30361;
wire n_30362;
wire n_30363;
wire n_30364;
wire n_30365;
wire n_30366;
wire n_30367;
wire n_30368;
wire n_30369;
wire n_30370;
wire n_30371;
wire n_30372;
wire n_30373;
wire n_30374;
wire n_30375;
wire n_30376;
wire n_30377;
wire n_30378;
wire n_30379;
wire n_30380;
wire n_30381;
wire n_30382;
wire n_30383;
wire n_30384;
wire n_30385;
wire n_30386;
wire n_30387;
wire n_30388;
wire n_30389;
wire n_30390;
wire n_30391;
wire n_30392;
wire n_30393;
wire n_30394;
wire n_30395;
wire n_30396;
wire n_30397;
wire n_30398;
wire n_30399;
wire n_30400;
wire n_30401;
wire n_30402;
wire n_30403;
wire n_30404;
wire n_30405;
wire n_30406;
wire n_30407;
wire n_30408;
wire n_30409;
wire n_30410;
wire n_30411;
wire n_30412;
wire n_30413;
wire n_30414;
wire n_30415;
wire n_30416;
wire n_30417;
wire n_30418;
wire n_30419;
wire n_30420;
wire n_30421;
wire n_30422;
wire n_30423;
wire n_30424;
wire n_30425;
wire n_30426;
wire n_30427;
wire n_30428;
wire n_30429;
wire n_30430;
wire n_30431;
wire n_30432;
wire n_30433;
wire n_30434;
wire n_30435;
wire n_30436;
wire n_30437;
wire n_30438;
wire n_30439;
wire n_30440;
wire n_30441;
wire n_30442;
wire n_30443;
wire n_30444;
wire n_30445;
wire n_30446;
wire n_30447;
wire n_30448;
wire n_30449;
wire n_30450;
wire n_30451;
wire n_30452;
wire n_30453;
wire n_30454;
wire n_30455;
wire n_30456;
wire n_30457;
wire n_30458;
wire n_30459;
wire n_30460;
wire n_30461;
wire n_30462;
wire n_30463;
wire n_30464;
wire n_30465;
wire n_30466;
wire n_30467;
wire n_30468;
wire n_30469;
wire n_30470;
wire n_30471;
wire n_30472;
wire n_30473;
wire n_30474;
wire n_30475;
wire n_30476;
wire n_30477;
wire n_30478;
wire n_30479;
wire n_30480;
wire n_30481;
wire n_30482;
wire n_30483;
wire n_30484;
wire n_30485;
wire n_30486;
wire n_30487;
wire n_30488;
wire n_30489;
wire n_30490;
wire n_30491;
wire n_30492;
wire n_30493;
wire n_30494;
wire n_30495;
wire n_30496;
wire n_30497;
wire n_30498;
wire n_30499;
wire n_30500;
wire n_30501;
wire n_30502;
wire n_30503;
wire n_30504;
wire n_30505;
wire n_30506;
wire n_30507;
wire n_30508;
wire n_30509;
wire n_30510;
wire n_30511;
wire n_30512;
wire n_30513;
wire n_30514;
wire n_30515;
wire n_30516;
wire n_30517;
wire n_30518;
wire n_30519;
wire n_30520;
wire n_30521;
wire n_30522;
wire n_30523;
wire n_30524;
wire n_30525;
wire n_30526;
wire n_30527;
wire n_30528;
wire n_30529;
wire n_30530;
wire n_30531;
wire n_30532;
wire n_30533;
wire n_30534;
wire n_30535;
wire n_30536;
wire n_30537;
wire n_30538;
wire n_30539;
wire n_30540;
wire n_30541;
wire n_30542;
wire n_30543;
wire n_30544;
wire n_30545;
wire n_30546;
wire n_30547;
wire n_30548;
wire n_30549;
wire n_30550;
wire n_30551;
wire n_30552;
wire n_30553;
wire n_30554;
wire n_30555;
wire n_30556;
wire n_30557;
wire n_30558;
wire n_30559;
wire n_30560;
wire n_30561;
wire n_30562;
wire n_30563;
wire n_30564;
wire n_30565;
wire n_30566;
wire n_30567;
wire n_30568;
wire n_30569;
wire n_30570;
wire n_30571;
wire n_30572;
wire n_30573;
wire n_30574;
wire n_30575;
wire n_30576;
wire n_30577;
wire n_30578;
wire n_30579;
wire n_30580;
wire n_30581;
wire n_30582;
wire n_30583;
wire n_30584;
wire n_30585;
wire n_30586;
wire n_30587;
wire n_30588;
wire n_30589;
wire n_30590;
wire n_30591;
wire n_30592;
wire n_30593;
wire n_30594;
wire n_30595;
wire n_30596;
wire n_30597;
wire n_30598;
wire n_30599;
wire n_30600;
wire n_30601;
wire n_30602;
wire n_30603;
wire n_30604;
wire n_30605;
wire n_30606;
wire n_30607;
wire n_30608;
wire n_30609;
wire n_30610;
wire n_30611;
wire n_30612;
wire n_30613;
wire n_30614;
wire n_30615;
wire n_30616;
wire n_30617;
wire n_30618;
wire n_30619;
wire n_30620;
wire n_30621;
wire n_30622;
wire n_30623;
wire n_30624;
wire n_30625;
wire n_30626;
wire n_30627;
wire n_30628;
wire n_30629;
wire n_30630;
wire n_30631;
wire n_30632;
wire n_30633;
wire n_30634;
wire n_30635;
wire n_30636;
wire n_30637;
wire n_30638;
wire n_30639;
wire n_30640;
wire n_30641;
wire n_30642;
wire n_30643;
wire n_30644;
wire n_30645;
wire n_30646;
wire n_30647;
wire n_30648;
wire n_30649;
wire n_30650;
wire n_30651;
wire n_30652;
wire n_30653;
wire n_30654;
wire n_30655;
wire n_30656;
wire n_30657;
wire n_30658;
wire n_30659;
wire n_30660;
wire n_30661;
wire n_30662;
wire n_30663;
wire n_30664;
wire n_30665;
wire n_30666;
wire n_30667;
wire n_30668;
wire n_30669;
wire n_30670;
wire n_30671;
wire n_30672;
wire n_30673;
wire n_30674;
wire n_30675;
wire n_30676;
wire n_30677;
wire n_30678;
wire n_30679;
wire n_30680;
wire n_30681;
wire n_30682;
wire n_30683;
wire n_30684;
wire n_30685;
wire n_30686;
wire n_30687;
wire n_30688;
wire n_30689;
wire n_30690;
wire n_30691;
wire n_30692;
wire n_30693;
wire n_30694;
wire n_30695;
wire n_30696;
wire n_30697;
wire n_30698;
wire n_30699;
wire n_30700;
wire n_30701;
wire n_30702;
wire n_30703;
wire n_30704;
wire n_30705;
wire n_30706;
wire n_30707;
wire n_30708;
wire n_30709;
wire n_30710;
wire n_30711;
wire n_30712;
wire n_30713;
wire n_30714;
wire n_30715;
wire n_30716;
wire n_30717;
wire n_30718;
wire n_30719;
wire n_30720;
wire n_30721;
wire n_30722;
wire n_30723;
wire n_30724;
wire n_30725;
wire n_30726;
wire n_30727;
wire n_30728;
wire n_30729;
wire n_30730;
wire n_30731;
wire n_30732;
wire n_30733;
wire n_30734;
wire n_30735;
wire n_30736;
wire n_30737;
wire n_30738;
wire n_30739;
wire n_30740;
wire n_30741;
wire n_30742;
wire n_30743;
wire n_30744;
wire n_30745;
wire n_30746;
wire n_30747;
wire n_30748;
wire n_30749;
wire n_30750;
wire n_30751;
wire n_30752;
wire n_30753;
wire n_30754;
wire n_30755;
wire n_30756;
wire n_30757;
wire n_30758;
wire n_30759;
wire n_30760;
wire n_30761;
wire n_30762;
wire n_30763;
wire n_30764;
wire n_30765;
wire n_30766;
wire n_30767;
wire n_30768;
wire n_30769;
wire n_30770;
wire n_30771;
wire n_30772;
wire n_30773;
wire n_30774;
wire n_30775;
wire n_30776;
wire n_30777;
wire n_30778;
wire n_30779;
wire n_30780;
wire n_30781;
wire n_30782;
wire n_30783;
wire n_30784;
wire n_30785;
wire n_30786;
wire n_30787;
wire n_30788;
wire n_30789;
wire n_30790;
wire n_30791;
wire n_30792;
wire n_30793;
wire n_30794;
wire n_30795;
wire n_30796;
wire n_30797;
wire n_30798;
wire n_30799;
wire n_30800;
wire n_30801;
wire n_30802;
wire n_30803;
wire n_30804;
wire n_30805;
wire n_30806;
wire n_30807;
wire n_30808;
wire n_30809;
wire n_30810;
wire n_30811;
wire n_30812;
wire n_30813;
wire n_30814;
wire n_30815;
wire n_30816;
wire n_30817;
wire n_30818;
wire n_30819;
wire n_30820;
wire n_30821;
wire n_30822;
wire n_30823;
wire n_30824;
wire n_30825;
wire n_30826;
wire n_30827;
wire n_30828;
wire n_30829;
wire n_30830;
wire n_30831;
wire n_30832;
wire n_30833;
wire n_30834;
wire n_30835;
wire n_30836;
wire n_30837;
wire n_30838;
wire n_30839;
wire n_30840;
wire n_30841;
wire n_30842;
wire n_30843;
wire n_30844;
wire n_30845;
wire n_30846;
wire n_30847;
wire n_30848;
wire n_30849;
wire n_30850;
wire n_30851;
wire n_30852;
wire n_30853;
wire n_30854;
wire n_30855;
wire n_30856;
wire n_30857;
wire n_30858;
wire n_30859;
wire n_30860;
wire n_30861;
wire n_30862;
wire n_30863;
wire n_30864;
wire n_30865;
wire n_30866;
wire n_30867;
wire n_30868;
wire n_30869;
wire n_30870;
wire n_30871;
wire n_30872;
wire n_30873;
wire n_30874;
wire n_30875;
wire n_30876;
wire n_30877;
wire n_30878;
wire n_30879;
wire n_30880;
wire n_30881;
wire n_30882;
wire n_30883;
wire n_30884;
wire n_30885;
wire n_30886;
wire n_30887;
wire n_30888;
wire n_30889;
wire n_30890;
wire n_30891;
wire n_30892;
wire n_30893;
wire n_30894;
wire n_30895;
wire n_30896;
wire n_30897;
wire n_30898;
wire n_30899;
wire n_30900;
wire n_30901;
wire n_30902;
wire n_30903;
wire n_30904;
wire n_30905;
wire n_30906;
wire n_30907;
wire n_30908;
wire n_30909;
wire n_30910;
wire n_30911;
wire n_30912;
wire n_30913;
wire n_30914;
wire n_30915;
wire n_30916;
wire n_30917;
wire n_30918;
wire n_30919;
wire n_30920;
wire n_30921;
wire n_30922;
wire n_30923;
wire n_30924;
wire n_30925;
wire n_30926;
wire n_30927;
wire n_30928;
wire n_30929;
wire n_30930;
wire n_30931;
wire n_30932;
wire n_30933;
wire n_30934;
wire n_30935;
wire n_30936;
wire n_30937;
wire n_30938;
wire n_30939;
wire n_30940;
wire n_30941;
wire n_30942;
wire n_30943;
wire n_30944;
wire n_30945;
wire n_30946;
wire n_30947;
wire n_30948;
wire n_30949;
wire n_30950;
wire n_30951;
wire n_30952;
wire n_30953;
wire n_30954;
wire n_30955;
wire n_30956;
wire n_30957;
wire n_30958;
wire n_30959;
wire n_30960;
wire n_30961;
wire n_30962;
wire n_30963;
wire n_30964;
wire n_30965;
wire n_30966;
wire n_30967;
wire n_30968;
wire n_30969;
wire n_30970;
wire n_30971;
wire n_30972;
wire n_30973;
wire n_30974;
wire n_30975;
wire n_30976;
wire n_30977;
wire n_30978;
wire n_30979;
wire n_30980;
wire n_30981;
wire n_30982;
wire n_30983;
wire n_30984;
wire n_30985;
wire n_30986;
wire n_30987;
wire n_30988;
wire n_30989;
wire n_30990;
wire n_30991;
wire n_30992;
wire n_30993;
wire n_30994;
wire n_30995;
wire n_30996;
wire n_30997;
wire n_30998;
wire n_30999;
wire n_31000;
wire n_31001;
wire n_31002;
wire n_31003;
wire n_31004;
wire n_31005;
wire n_31006;
wire n_31007;
wire n_31008;
wire n_31009;
wire n_31010;
wire n_31011;
wire n_31012;
wire n_31013;
wire n_31014;
wire n_31015;
wire n_31016;
wire n_31017;
wire n_31018;
wire n_31019;
wire n_31020;
wire n_31021;
wire n_31022;
wire n_31023;
wire n_31024;
wire n_31025;
wire n_31026;
wire n_31027;
wire n_31028;
wire n_31029;
wire n_31030;
wire n_31031;
wire n_31032;
wire n_31033;
wire n_31034;
wire n_31035;
wire n_31036;
wire n_31037;
wire n_31038;
wire n_31039;
wire n_31040;
wire n_31041;
wire n_31042;
wire n_31043;
wire n_31044;
wire n_31045;
wire n_31046;
wire n_31047;
wire n_31048;
wire n_31049;
wire n_31050;
wire n_31051;
wire n_31052;
wire n_31053;
wire n_31054;
wire n_31055;
wire n_31056;
wire n_31057;
wire n_31058;
wire n_31059;
wire n_31060;
wire n_31061;
wire n_31062;
wire n_31063;
wire n_31064;
wire n_31065;
wire n_31066;
wire n_31067;
wire n_31068;
wire n_31069;
wire n_31070;
wire n_31071;
wire n_31072;
wire n_31073;
wire n_31074;
wire n_31075;
wire n_31076;
wire n_31077;
wire n_31078;
wire n_31079;
wire n_31080;
wire n_31081;
wire n_31082;
wire n_31083;
wire n_31084;
wire n_31085;
wire n_31086;
wire n_31087;
wire n_31088;
wire n_31089;
wire n_31090;
wire n_31091;
wire n_31092;
wire n_31093;
wire n_31094;
wire n_31095;
wire n_31096;
wire n_31097;
wire n_31098;
wire n_31099;
wire n_31100;
wire n_31101;
wire n_31102;
wire n_31103;
wire n_31104;
wire n_31105;
wire n_31106;
wire n_31107;
wire n_31108;
wire n_31109;
wire n_31110;
wire n_31111;
wire n_31112;
wire n_31113;
wire n_31114;
wire n_31115;
wire n_31116;
wire n_31117;
wire n_31118;
wire n_31119;
wire n_31120;
wire n_31121;
wire n_31122;
wire n_31123;
wire n_31124;
wire n_31125;
wire n_31126;
wire n_31127;
wire n_31128;
wire n_31129;
wire n_31130;
wire n_31131;
wire n_31132;
wire n_31133;
wire n_31134;
wire n_31135;
wire n_31136;
wire n_31137;
wire n_31138;
wire n_31139;
wire n_31140;
wire n_31141;
wire n_31142;
wire n_31143;
wire n_31144;
wire n_31145;
wire n_31146;
wire n_31147;
wire n_31148;
wire n_31149;
wire n_31150;
wire n_31151;
wire n_31152;
wire n_31153;
wire n_31154;
wire n_31155;
wire n_31156;
wire n_31157;
wire n_31158;
wire n_31159;
wire n_31160;
wire n_31161;
wire n_31162;
wire n_31163;
wire n_31164;
wire n_31165;
wire n_31166;
wire n_31167;
wire n_31168;
wire n_31169;
wire n_31170;
wire n_31171;
wire n_31172;
wire n_31173;
wire n_31174;
wire n_31175;
wire n_31176;
wire n_31177;
wire n_31178;
wire n_31179;
wire n_31180;
wire n_31181;
wire n_31182;
wire n_31183;
wire n_31184;
wire n_31185;
wire n_31186;
wire n_31187;
wire n_31188;
wire n_31189;
wire n_31190;
wire n_31191;
wire n_31192;
wire n_31193;
wire n_31194;
wire n_31195;
wire n_31196;
wire n_31197;
wire n_31198;
wire n_31199;
wire n_31200;
wire n_31201;
wire n_31202;
wire n_31203;
wire n_31204;
wire n_31205;
wire n_31206;
wire n_31207;
wire n_31208;
wire n_31209;
wire n_31210;
wire n_31211;
wire n_31212;
wire n_31213;
wire n_31214;
wire n_31215;
wire n_31216;
wire n_31217;
wire n_31218;
wire n_31219;
wire n_31220;
wire n_31221;
wire n_31222;
wire n_31223;
wire n_31224;
wire n_31225;
wire n_31226;
wire n_31227;
wire n_31228;
wire n_31229;
wire n_31230;
wire n_31231;
wire n_31232;
wire n_31233;
wire n_31234;
wire n_31235;
wire n_31236;
wire n_31237;
wire n_31238;
wire n_31239;
wire n_31240;
wire n_31241;
wire n_31242;
wire n_31243;
wire n_31244;
wire n_31245;
wire n_31246;
wire n_31247;
wire n_31248;
wire n_31249;
wire n_31250;
wire n_31251;
wire n_31252;
wire n_31253;
wire n_31254;
wire n_31255;
wire n_31256;
wire n_31257;
wire n_31258;
wire n_31259;
wire n_31260;
wire n_31261;
wire n_31262;
wire n_31263;
wire n_31264;
wire n_31265;
wire n_31266;
wire n_31267;
wire n_31268;
wire n_31269;
wire n_31270;
wire n_31271;
wire n_31272;
wire n_31273;
wire n_31274;
wire n_31275;
wire n_31276;
wire n_31277;
wire n_31278;
wire n_31279;
wire n_31280;
wire n_31281;
wire n_31282;
wire n_31283;
wire n_31284;
wire n_31285;
wire n_31286;
wire n_31287;
wire n_31288;
wire n_31289;
wire n_31290;
wire n_31291;
wire n_31292;
wire n_31293;
wire n_31294;
wire n_31295;
wire n_31296;
wire n_31297;
wire n_31298;
wire n_31299;
wire n_31300;
wire n_31301;
wire n_31302;
wire n_31303;
wire n_31304;
wire n_31305;
wire n_31306;
wire n_31307;
wire n_31308;
wire n_31309;
wire n_31310;
wire n_31311;
wire n_31312;
wire n_31313;
wire n_31314;
wire n_31315;
wire n_31316;
wire n_31317;
wire n_31318;
wire n_31319;
wire n_31320;
wire n_31321;
wire n_31322;
wire n_31323;
wire n_31324;
wire n_31325;
wire n_31326;
wire n_31327;
wire n_31328;
wire n_31329;
wire n_31330;
wire n_31331;
wire n_31332;
wire n_31333;
wire n_31334;
wire n_31335;
wire n_31336;
wire n_31337;
wire n_31338;
wire n_31339;
wire n_31340;
wire n_31341;
wire n_31342;
wire n_31343;
wire n_31344;
wire n_31345;
wire n_31346;
wire n_31347;
wire n_31348;
wire n_31349;
wire n_31350;
wire n_31351;
wire n_31352;
wire n_31353;
wire n_31354;
wire n_31355;
wire n_31356;
wire n_31357;
wire n_31358;
wire n_31359;
wire n_31360;
wire n_31361;
wire n_31362;
wire n_31363;
wire n_31364;
wire n_31365;
wire n_31366;
wire n_31367;
wire n_31368;
wire n_31369;
wire n_31370;
wire n_31371;
wire n_31372;
wire n_31373;
wire n_31374;
wire n_31375;
wire n_31376;
wire n_31377;
wire n_31378;
wire n_31379;
wire n_31380;
wire n_31381;
wire n_31382;
wire n_31383;
wire n_31384;
wire n_31385;
wire n_31386;
wire n_31387;
wire n_31388;
wire n_31389;
wire n_31390;
wire n_31391;
wire n_31392;
wire n_31393;
wire n_31394;
wire n_31395;
wire n_31396;
wire n_31397;
wire n_31398;
wire n_31399;
wire n_31400;
wire n_31401;
wire n_31402;
wire n_31403;
wire n_31404;
wire n_31405;
wire n_31406;
wire n_31407;
wire n_31408;
wire n_31409;
wire n_31410;
wire n_31411;
wire n_31412;
wire n_31413;
wire n_31414;
wire n_31415;
wire n_31416;
wire n_31417;
wire n_31418;
wire n_31419;
wire n_31420;
wire n_31421;
wire n_31422;
wire n_31423;
wire n_31424;
wire n_31425;
wire n_31426;
wire n_31427;
wire n_31428;
wire n_31429;
wire n_31430;
wire n_31431;
wire n_31432;
wire n_31433;
wire n_31434;
wire n_31435;
wire n_31436;
wire n_31437;
wire n_31438;
wire n_31439;
wire n_31440;
wire n_31441;
wire n_31442;
wire n_31443;
wire n_31444;
wire n_31445;
wire n_31446;
wire n_31447;
wire n_31448;
wire n_31449;
wire n_31450;
wire n_31451;
wire n_31452;
wire n_31453;
wire n_31454;
wire n_31455;
wire n_31456;
wire n_31457;
wire n_31458;
wire n_31459;
wire n_31460;
wire n_31461;
wire n_31462;
wire n_31463;
wire n_31464;
wire n_31465;
wire n_31466;
wire n_31467;
wire n_31468;
wire n_31469;
wire n_31470;
wire n_31471;
wire n_31472;
wire n_31473;
wire n_31474;
wire n_31475;
wire n_31476;
wire n_31477;
wire n_31478;
wire n_31479;
wire n_31480;
wire n_31481;
wire n_31482;
wire n_31483;
wire n_31484;
wire n_31485;
wire n_31486;
wire n_31487;
wire n_31488;
wire n_31489;
wire n_31490;
wire n_31491;
wire n_31492;
wire n_31493;
wire n_31494;
wire n_31495;
wire n_31496;
wire n_31497;
wire n_31498;
wire n_31499;
wire n_31500;
wire n_31501;
wire n_31502;
wire n_31503;
wire n_31504;
wire n_31505;
wire n_31506;
wire n_31507;
wire n_31508;
wire n_31509;
wire n_31510;
wire n_31511;
wire n_31512;
wire n_31513;
wire n_31514;
wire n_31515;
wire n_31516;
wire n_31517;
wire n_31518;
wire n_31519;
wire n_31520;
wire n_31521;
wire n_31522;
wire n_31523;
wire n_31524;
wire n_31525;
wire n_31526;
wire n_31527;
wire n_31528;
wire n_31529;
wire n_31530;
wire n_31531;
wire n_31532;
wire n_31533;
wire n_31534;
wire n_31535;
wire n_31536;
wire n_31537;
wire n_31538;
wire n_31539;
wire n_31540;
wire n_31541;
wire n_31542;
wire n_31543;
wire n_31544;
wire n_31545;
wire n_31546;
wire n_31547;
wire n_31548;
wire n_31549;
wire n_31550;
wire n_31551;
wire n_31552;
wire n_31553;
wire n_31554;
wire n_31555;
wire n_31556;
wire n_31557;
wire n_31558;
wire n_31559;
wire n_31560;
wire n_31561;
wire n_31562;
wire n_31563;
wire n_31564;
wire n_31565;
wire n_31566;
wire n_31567;
wire n_31568;
wire n_31569;
wire n_31570;
wire n_31571;
wire n_31572;
wire n_31573;
wire n_31574;
wire n_31575;
wire n_31576;
wire n_31577;
wire n_31578;
wire n_31579;
wire n_31580;
wire n_31581;
wire n_31582;
wire n_31583;
wire n_31584;
wire n_31585;
wire n_31586;
wire n_31587;
wire n_31588;
wire n_31589;
wire n_31590;
wire n_31591;
wire n_31592;
wire n_31593;
wire n_31594;
wire n_31595;
wire n_31596;
wire n_31597;
wire n_31598;
wire n_31599;
wire n_31600;
wire n_31601;
wire n_31602;
wire n_31603;
wire n_31604;
wire n_31605;
wire n_31606;
wire n_31607;
wire n_31608;
wire n_31609;
wire n_31610;
wire n_31611;
wire n_31612;
wire n_31613;
wire n_31614;
wire n_31615;
wire n_31616;
wire n_31617;
wire n_31618;
wire n_31619;
wire n_31620;
wire n_31621;
wire n_31622;
wire n_31623;
wire n_31624;
wire n_31625;
wire n_31626;
wire n_31627;
wire n_31628;
wire n_31629;
wire n_31630;
wire n_31631;
wire n_31632;
wire n_31633;
wire n_31634;
wire n_31635;
wire n_31636;
wire n_31637;
wire n_31638;
wire n_31639;
wire n_31640;
wire n_31641;
wire n_31642;
wire n_31643;
wire n_31644;
wire n_31645;
wire n_31646;
wire n_31647;
wire n_31648;
wire n_31649;
wire n_31650;
wire n_31651;
wire n_31652;
wire n_31653;
wire n_31654;
wire n_31655;
wire n_31656;
wire n_31657;
wire n_31658;
wire n_31659;
wire n_31660;
wire n_31661;
wire n_31662;
wire n_31663;
wire n_31664;
wire n_31665;
wire n_31666;
wire n_31667;
wire n_31668;
wire n_31669;
wire n_31670;
wire n_31671;
wire n_31672;
wire n_31673;
wire n_31674;
wire n_31675;
wire n_31676;
wire n_31677;
wire n_31678;
wire n_31679;
wire n_31680;
wire n_31681;
wire n_31682;
wire n_31683;
wire n_31684;
wire n_31685;
wire n_31686;
wire n_31687;
wire n_31688;
wire n_31689;
wire n_31690;
wire n_31691;
wire n_31692;
wire n_31693;
wire n_31694;
wire n_31695;
wire n_31696;
wire n_31697;
wire n_31698;
wire n_31699;
wire n_31700;
wire n_31701;
wire n_31702;
wire n_31703;
wire n_31704;
wire n_31705;
wire n_31706;
wire n_31707;
wire n_31708;
wire n_31709;
wire n_31710;
wire n_31711;
wire n_31712;
wire n_31713;
wire n_31714;
wire n_31715;
wire n_31716;
wire n_31717;
wire n_31718;
wire n_31719;
wire n_31720;
wire n_31721;
wire n_31722;
wire n_31723;
wire n_31724;
wire n_31725;
wire n_31726;
wire n_31727;
wire n_31728;
wire n_31729;
wire n_31730;
wire n_31731;
wire n_31732;
wire n_31733;
wire n_31734;
wire n_31735;
wire n_31736;
wire n_31737;
wire n_31738;
wire n_31739;
wire n_31740;
wire n_31741;
wire n_31742;
wire n_31743;
wire n_31744;
wire n_31745;
wire n_31746;
wire n_31747;
wire n_31748;
wire n_31749;
wire n_31750;
wire n_31751;
wire n_31752;
wire n_31753;
wire n_31754;
wire n_31755;
wire n_31756;
wire n_31757;
wire n_31758;
wire n_31759;
wire n_31760;
wire n_31761;
wire n_31762;
wire n_31763;
wire n_31764;
wire n_31765;
wire n_31766;
wire n_31767;
wire n_31768;
wire n_31769;
wire n_31770;
wire n_31771;
wire n_31772;
wire n_31773;
wire n_31774;
wire n_31775;
wire n_31776;
wire n_31777;
wire n_31778;
wire n_31779;
wire n_31780;
wire n_31781;
wire n_31782;
wire n_31783;
wire n_31784;
wire n_31785;
wire n_31786;
wire n_31787;
wire n_31788;
wire n_31789;
wire n_31790;
wire n_31791;
wire n_31792;
wire n_31793;
wire n_31794;
wire n_31795;
wire n_31796;
wire n_31797;
wire n_31798;
wire n_31799;
wire n_31800;
wire n_31801;
wire n_31802;
wire n_31803;
wire n_31804;
wire n_31805;
wire n_31806;
wire n_31807;
wire n_31808;
wire n_31809;
wire n_31810;
wire n_31811;
wire n_31812;
wire n_31813;
wire n_31814;
wire n_31815;
wire n_31816;
wire n_31817;
wire n_31818;
wire n_31819;
wire n_31820;
wire n_31821;
wire n_31822;
wire n_31823;
wire n_31824;
wire n_31825;
wire n_31826;
wire n_31827;
wire n_31828;
wire n_31829;
wire n_31830;
wire n_31831;
wire n_31832;
wire n_31833;
wire n_31834;
wire n_31835;
wire n_31836;
wire n_31837;
wire n_31838;
wire n_31839;
wire n_31840;
wire n_31841;
wire n_31842;
wire n_31843;
wire n_31844;
wire n_31845;
wire n_31846;
wire n_31847;
wire n_31848;
wire n_31849;
wire n_31850;
wire n_31851;
wire n_31852;
wire n_31853;
wire n_31854;
wire n_31855;
wire n_31856;
wire n_31857;
wire n_31858;
wire n_31859;
wire n_31860;
wire n_31861;
wire n_31862;
wire n_31863;
wire n_31864;
wire n_31865;
wire n_31866;
wire n_31867;
wire n_31868;
wire n_31869;
wire n_31870;
wire n_31871;
wire n_31872;
wire n_31873;
wire n_31874;
wire n_31875;
wire n_31876;
wire n_31877;
wire n_31878;
wire n_31879;
wire n_31880;
wire n_31881;
wire n_31882;
wire n_31883;
wire n_31884;
wire n_31885;
wire n_31886;
wire n_31887;
wire n_31888;
wire n_31889;
wire n_31890;
wire n_31891;
wire n_31892;
wire n_31893;
wire n_31894;
wire n_31895;
wire n_31896;
wire n_31897;
wire n_31898;
wire n_31899;
wire n_31900;
wire n_31901;
wire n_31902;
wire n_31903;
wire n_31904;
wire n_31905;
wire n_31906;
wire n_31907;
wire n_31908;
wire n_31909;
wire n_31910;
wire n_31911;
wire n_31912;
wire n_31913;
wire n_31914;
wire n_31915;
wire n_31916;
wire n_31917;
wire n_31918;
wire n_31919;
wire n_31920;
wire n_31921;
wire n_31922;
wire n_31923;
wire n_31924;
wire n_31925;
wire n_31926;
wire n_31927;
wire n_31928;
wire n_31929;
wire n_31930;
wire n_31931;
wire n_31932;
wire n_31933;
wire n_31934;
wire n_31935;
wire n_31936;
wire n_31937;
wire n_31938;
wire n_31939;
wire n_31940;
wire n_31941;
wire n_31942;
wire n_31943;
wire n_31944;
wire n_31945;
wire n_31946;
wire n_31947;
wire n_31948;
wire n_31949;
wire n_31950;
wire n_31951;
wire n_31952;
wire n_31953;
wire n_31954;
wire n_31955;
wire n_31956;
wire n_31957;
wire n_31958;
wire n_31959;
wire n_31960;
wire n_31961;
wire n_31962;
wire n_31963;
wire n_31964;
wire n_31965;
wire n_31966;
wire n_31967;
wire n_31968;
wire n_31969;
wire n_31970;
wire n_31971;
wire n_31972;
wire n_31973;
wire n_31974;
wire n_31975;
wire n_31976;
wire n_31977;
wire n_31978;
wire n_31979;
wire n_31980;
wire n_31981;
wire n_31982;
wire n_31983;
wire n_31984;
wire n_31985;
wire n_31986;
wire n_31987;
wire n_31988;
wire n_31989;
wire n_31990;
wire n_31991;
wire n_31992;
wire n_31993;
wire n_31994;
wire n_31995;
wire n_31996;
wire n_31997;
wire n_31998;
wire n_31999;
wire n_32000;
wire n_32001;
wire n_32002;
wire n_32003;
wire n_32004;
wire n_32005;
wire n_32006;
wire n_32007;
wire n_32008;
wire n_32009;
wire n_32010;
wire n_32011;
wire n_32012;
wire n_32013;
wire n_32014;
wire n_32015;
wire n_32016;
wire n_32017;
wire n_32018;
wire n_32019;
wire n_32020;
wire n_32021;
wire n_32022;
wire n_32023;
wire n_32024;
wire n_32025;
wire n_32026;
wire n_32027;
wire n_32028;
wire n_32029;
wire n_32030;
wire n_32031;
wire n_32032;
wire n_32033;
wire n_32034;
wire n_32035;
wire n_32036;
wire n_32037;
wire n_32038;
wire n_32039;
wire n_32040;
wire n_32041;
wire n_32042;
wire n_32043;
wire n_32044;
wire n_32045;
wire n_32046;
wire n_32047;
wire n_32048;
wire n_32049;
wire n_32050;
wire n_32051;
wire n_32052;
wire n_32053;
wire n_32054;
wire n_32055;
wire n_32056;
wire n_32057;
wire n_32058;
wire n_32059;
wire n_32060;
wire n_32061;
wire n_32062;
wire n_32063;
wire n_32064;
wire n_32065;
wire n_32066;
wire n_32067;
wire n_32068;
wire n_32069;
wire n_32070;
wire n_32071;
wire n_32072;
wire n_32073;
wire n_32074;
wire n_32075;
wire n_32076;
wire n_32077;
wire n_32078;
wire n_32079;
wire n_32080;
wire n_32081;
wire n_32082;
wire n_32083;
wire n_32084;
wire n_32085;
wire n_32086;
wire n_32087;
wire n_32088;
wire n_32089;
wire n_32090;
wire n_32091;
wire n_32092;
wire n_32093;
wire n_32094;
wire n_32095;
wire n_32096;
wire n_32097;
wire n_32098;
wire n_32099;
wire n_32100;
wire n_32101;
wire n_32102;
wire n_32103;
wire n_32104;
wire n_32105;
wire n_32106;
wire n_32107;
wire n_32108;
wire n_32109;
wire n_32110;
wire n_32111;
wire n_32112;
wire n_32113;
wire n_32114;
wire n_32115;
wire n_32116;
wire n_32117;
wire n_32118;
wire n_32119;
wire n_32120;
wire n_32121;
wire n_32122;
wire n_32123;
wire n_32124;
wire n_32125;
wire n_32126;
wire n_32127;
wire n_32128;
wire n_32129;
wire n_32130;
wire n_32131;
wire n_32132;
wire n_32133;
wire n_32134;
wire n_32135;
wire n_32136;
wire n_32137;
wire n_32138;
wire n_32139;
wire n_32140;
wire n_32141;
wire n_32142;
wire n_32143;
wire n_32144;
wire n_32145;
wire n_32146;
wire n_32147;
wire n_32148;
wire n_32149;
wire n_32150;
wire n_32151;
wire n_32152;
wire n_32153;
wire n_32154;
wire n_32155;
wire n_32156;
wire n_32157;
wire n_32158;
wire n_32159;
wire n_32160;
wire n_32161;
wire n_32162;
wire n_32163;
wire n_32164;
wire n_32165;
wire n_32166;
wire n_32167;
wire n_32168;
wire n_32169;
wire n_32170;
wire n_32171;
wire n_32172;
wire n_32173;
wire n_32174;
wire n_32175;
wire n_32176;
wire n_32177;
wire n_32178;
wire n_32179;
wire n_32180;
wire n_32181;
wire n_32182;
wire n_32183;
wire n_32184;
wire n_32185;
wire n_32186;
wire n_32187;
wire n_32188;
wire n_32189;
wire n_32190;
wire n_32191;
wire n_32192;
wire n_32193;
wire n_32194;
wire n_32195;
wire n_32196;
wire n_32197;
wire n_32198;
wire n_32199;
wire n_32200;
wire n_32201;
wire n_32202;
wire n_32203;
wire n_32204;
wire n_32205;
wire n_32206;
wire n_32207;
wire n_32208;
wire n_32209;
wire n_32210;
wire n_32211;
wire n_32212;
wire n_32213;
wire n_32214;
wire n_32215;
wire n_32216;
wire n_32217;
wire n_32218;
wire n_32219;
wire n_32220;
wire n_32221;
wire n_32222;
wire n_32223;
wire n_32224;
wire n_32225;
wire n_32226;
wire n_32227;
wire n_32228;
wire n_32229;
wire n_32230;
wire n_32231;
wire n_32232;
wire n_32233;
wire n_32234;
wire n_32235;
wire n_32236;
wire n_32237;
wire n_32238;
wire n_32239;
wire n_32240;
wire n_32241;
wire n_32242;
wire n_32243;
wire n_32244;
wire n_32245;
wire n_32246;
wire n_32247;
wire n_32248;
wire n_32249;
wire n_32250;
wire n_32251;
wire n_32252;
wire n_32253;
wire n_32254;
wire n_32255;
wire n_32256;
wire n_32257;
wire n_32258;
wire n_32259;
wire n_32260;
wire n_32261;
wire n_32262;
wire n_32263;
wire n_32264;
wire n_32265;
wire n_32266;
wire n_32267;
wire n_32268;
wire n_32269;
wire n_32270;
wire n_32271;
wire n_32272;
wire n_32273;
wire n_32274;
wire n_32275;
wire n_32276;
wire n_32277;
wire n_32278;
wire n_32279;
wire n_32280;
wire n_32281;
wire n_32282;
wire n_32283;
wire n_32284;
wire n_32285;
wire n_32286;
wire n_32287;
wire n_32288;
wire n_32289;
wire n_32290;
wire n_32291;
wire n_32292;
wire n_32293;
wire n_32294;
wire n_32295;
wire n_32296;
wire n_32297;
wire n_32298;
wire n_32299;
wire n_32300;
wire n_32301;
wire n_32302;
wire n_32303;
wire n_32304;
wire n_32305;
wire n_32306;
wire n_32307;
wire n_32308;
wire n_32309;
wire n_32310;
wire n_32311;
wire n_32312;
wire n_32313;
wire n_32314;
wire n_32315;
wire n_32316;
wire n_32317;
wire n_32318;
wire n_32319;
wire n_32320;
wire n_32321;
wire n_32322;
wire n_32323;
wire n_32324;
wire n_32325;
wire n_32326;
wire n_32327;
wire n_32328;
wire n_32329;
wire n_32330;
wire n_32331;
wire n_32332;
wire n_32333;
wire n_32334;
wire n_32335;
wire n_32336;
wire n_32337;
wire n_32338;
wire n_32339;
wire n_32340;
wire n_32341;
wire n_32342;
wire n_32343;
wire n_32344;
wire n_32345;
wire n_32346;
wire n_32347;
wire n_32348;
wire n_32349;
wire n_32350;
wire n_32351;
wire n_32352;
wire n_32353;
wire n_32354;
wire n_32355;
wire n_32356;
wire n_32357;
wire n_32358;
wire n_32359;
wire n_32360;
wire n_32361;
wire n_32362;
wire n_32363;
wire n_32364;
wire n_32365;
wire n_32366;
wire n_32367;
wire n_32368;
wire n_32369;
wire n_32370;
wire n_32371;
wire n_32372;
wire n_32373;
wire n_32374;
wire n_32375;
wire n_32376;
wire n_32377;
wire n_32378;
wire n_32379;
wire n_32380;
wire n_32381;
wire n_32382;
wire n_32383;
wire n_32384;
wire n_32385;
wire n_32386;
wire n_32387;
wire n_32388;
wire n_32389;
wire n_32390;
wire n_32391;
wire n_32392;
wire n_32393;
wire n_32394;
wire n_32395;
wire n_32396;
wire n_32397;
wire n_32398;
wire n_32399;
wire n_32400;
wire n_32401;
wire n_32402;
wire n_32403;
wire n_32404;
wire n_32405;
wire n_32406;
wire n_32407;
wire n_32408;
wire n_32409;
wire n_32410;
wire n_32411;
wire n_32412;
wire n_32413;
wire n_32414;
wire n_32415;
wire n_32416;
wire n_32417;
wire n_32418;
wire n_32419;
wire n_32420;
wire n_32421;
wire n_32422;
wire n_32423;
wire n_32424;
wire n_32425;
wire n_32426;
wire n_32427;
wire n_32428;
wire n_32429;
wire n_32430;
wire n_32431;
wire n_32432;
wire n_32433;
wire n_32434;
wire n_32435;
wire n_32436;
wire n_32437;
wire n_32438;
wire n_32439;
wire n_32440;
wire n_32441;
wire n_32442;
wire n_32443;
wire n_32444;
wire n_32445;
wire n_32446;
wire n_32447;
wire n_32448;
wire n_32449;
wire n_32450;
wire n_32451;
wire n_32452;
wire n_32453;
wire n_32454;
wire n_32455;
wire n_32456;
wire n_32457;
wire n_32458;
wire n_32459;
wire n_32460;
wire n_32461;
wire n_32462;
wire n_32463;
wire n_32464;
wire n_32465;
wire n_32466;
wire n_32467;
wire n_32468;
wire n_32469;
wire n_32470;
wire n_32471;
wire n_32472;
wire n_32473;
wire n_32474;
wire n_32475;
wire n_32476;
wire n_32477;
wire n_32478;
wire n_32479;
wire n_32480;
wire n_32481;
wire n_32482;
wire n_32483;
wire n_32484;
wire n_32485;
wire n_32486;
wire n_32487;
wire n_32488;
wire n_32489;
wire n_32490;
wire n_32491;
wire n_32492;
wire n_32493;
wire n_32494;
wire n_32495;
wire n_32496;
wire n_32497;
wire n_32498;
wire n_32499;
wire n_32500;
wire n_32501;
wire n_32502;
wire n_32503;
wire n_32504;
wire n_32505;
wire n_32506;
wire n_32507;
wire n_32508;
wire n_32509;
wire n_32510;
wire n_32511;
wire n_32512;
wire n_32513;
wire n_32514;
wire n_32515;
wire n_32516;
wire n_32517;
wire n_32518;
wire n_32519;
wire n_32520;
wire n_32521;
wire n_32522;
wire n_32523;
wire n_32524;
wire n_32525;
wire n_32526;
wire n_32527;
wire n_32528;
wire n_32529;
wire n_32530;
wire n_32531;
wire n_32532;
wire n_32533;
wire n_32534;
wire n_32535;
wire n_32536;
wire n_32537;
wire n_32538;
wire n_32539;
wire n_32540;
wire n_32541;
wire n_32542;
wire n_32543;
wire n_32544;
wire n_32545;
wire n_32546;
wire n_32547;
wire n_32548;
wire n_32549;
wire n_32550;
wire n_32551;
wire n_32552;
wire n_32553;
wire n_32554;
wire n_32555;
wire n_32556;
wire n_32557;
wire n_32558;
wire n_32559;
wire n_32560;
wire n_32561;
wire n_32562;
wire n_32563;
wire n_32564;
wire n_32565;
wire n_32566;
wire n_32567;
wire n_32568;
wire n_32569;
wire n_32570;
wire n_32571;
wire n_32572;
wire n_32573;
wire n_32574;
wire n_32575;
wire n_32576;
wire n_32577;
wire n_32578;
wire n_32579;
wire n_32580;
wire n_32581;
wire n_32582;
wire n_32583;
wire n_32584;
wire n_32585;
wire n_32586;
wire n_32587;
wire n_32588;
wire n_32589;
wire n_32590;
wire n_32591;
wire n_32592;
wire n_32593;
wire n_32594;
wire n_32595;
wire n_32596;
wire n_32597;
wire n_32598;
wire n_32599;
wire n_32600;
wire n_32601;
wire n_32602;
wire n_32603;
wire n_32604;
wire n_32605;
wire n_32606;
wire n_32607;
wire n_32608;
wire n_32609;
wire n_32610;
wire n_32611;
wire n_32612;
wire n_32613;
wire n_32614;
wire n_32615;
wire n_32616;
wire n_32617;
wire n_32618;
wire n_32619;
wire n_32620;
wire n_32621;
wire n_32622;
wire n_32623;
wire n_32624;
wire n_32625;
wire n_32626;
wire n_32627;
wire n_32628;
wire n_32629;
wire n_32630;
wire n_32631;
wire n_32632;
wire n_32633;
wire n_32634;
wire n_32635;
wire n_32636;
wire n_32637;
wire n_32638;
wire n_32639;
wire n_32640;
wire n_32641;
wire n_32642;
wire n_32643;
wire n_32644;
wire n_32645;
wire n_32646;
wire n_32647;
wire n_32648;
wire n_32649;
wire n_32650;
wire n_32651;
wire n_32652;
wire n_32653;
wire n_32654;
wire n_32655;
wire n_32656;
wire n_32657;
wire n_32658;
wire n_32659;
wire n_32660;
wire n_32661;
wire n_32662;
wire n_32663;
wire n_32664;
wire n_32665;
wire n_32666;
wire n_32667;
wire n_32668;
wire n_32669;
wire n_32670;
wire n_32671;
wire n_32672;
wire n_32673;
wire n_32674;
wire n_32675;
wire n_32676;
wire n_32677;
wire n_32678;
wire n_32679;
wire n_32680;
wire n_32681;
wire n_32682;
wire n_32683;
wire n_32684;
wire n_32685;
wire n_32686;
wire n_32687;
wire n_32688;
wire n_32689;
wire n_32690;
wire n_32691;
wire n_32692;
wire n_32693;
wire n_32694;
wire n_32695;
wire n_32696;
wire n_32697;
wire n_32698;
wire n_32699;
wire n_32700;
wire n_32701;
wire n_32702;
wire n_32703;
wire n_32704;
wire n_32705;
wire n_32706;
wire n_32707;
wire n_32708;
wire n_32709;
wire n_32710;
wire n_32711;
wire n_32712;
wire n_32713;
wire n_32714;
wire n_32715;
wire n_32716;
wire n_32717;
wire n_32718;
wire n_32719;
wire n_32720;
wire n_32721;
wire n_32722;
wire n_32723;
wire n_32724;
wire n_32725;
wire n_32726;
wire n_32727;
wire n_32728;
wire n_32729;
wire n_32730;
wire n_32731;
wire n_32732;
wire n_32733;
wire n_32734;
wire n_32735;
wire n_32736;
wire n_32737;
wire n_32738;
wire n_32739;
wire n_32740;
wire n_32741;
wire n_32742;
wire n_32743;
wire n_32744;
wire n_32745;
wire n_32746;
wire n_32747;
wire n_32748;
wire n_32749;
wire n_32750;
wire n_32751;
wire n_32752;
wire n_32753;
wire n_32754;
wire n_32755;
wire n_32756;
wire n_32757;
wire n_32758;
wire n_32759;
wire n_32760;
wire n_32761;
wire n_32762;
wire n_32763;
wire n_32764;
wire n_32765;
wire n_32766;
wire n_32767;
wire n_32768;
wire n_32769;
wire n_32770;
wire n_32771;
wire n_32772;
wire n_32773;
wire n_32774;
wire n_32775;
wire n_32776;
wire n_32777;
wire n_32778;
wire n_32779;
wire n_32780;
wire n_32781;
wire n_32782;
wire n_32783;
wire n_32784;
wire n_32785;
wire n_32786;
wire n_32787;
wire n_32788;
wire n_32789;
wire n_32790;
wire n_32791;
wire n_32792;
wire n_32793;
wire n_32794;
wire n_32795;
wire n_32796;
wire n_32797;
wire n_32798;
wire n_32799;
wire n_32800;
wire n_32801;
wire n_32802;
wire n_32803;
wire n_32804;
wire n_32805;
wire n_32806;
wire n_32807;
wire n_32808;
wire n_32809;
wire n_32810;
wire n_32811;
wire n_32812;
wire n_32813;
wire n_32814;
wire n_32815;
wire n_32816;
wire n_32817;
wire n_32818;
wire n_32819;
wire n_32820;
wire n_32821;
wire n_32822;
wire n_32823;
wire n_32824;
wire n_32825;
wire n_32826;
wire n_32827;
wire n_32828;
wire n_32829;
wire n_32830;
wire n_32831;
wire n_32832;
wire n_32833;
wire n_32834;
wire n_32835;
wire n_32836;
wire n_32837;
wire n_32838;
wire n_32839;
wire n_32840;
wire n_32841;
wire n_32842;
wire n_32843;
wire n_32844;
wire n_32845;
wire n_32846;
wire n_32847;
wire n_32848;
wire n_32849;
wire n_32850;
wire n_32851;
wire n_32852;
wire n_32853;
wire n_32854;
wire n_32855;
wire n_32856;
wire n_32857;
wire n_32858;
wire n_32859;
wire n_32860;
wire n_32861;
wire n_32862;
wire n_32863;
wire n_32864;
wire n_32865;
wire n_32866;
wire n_32867;
wire n_32868;
wire n_32869;
wire n_32870;
wire n_32871;
wire n_32872;
wire n_32873;
wire n_32874;
wire n_32875;
wire n_32876;
wire n_32877;
wire n_32878;
wire n_32879;
wire n_32880;
wire n_32881;
wire n_32882;
wire n_32883;
wire n_32884;
wire n_32885;
wire n_32886;
wire n_32887;
wire n_32888;
wire n_32889;
wire n_32890;
wire n_32891;
wire n_32892;
wire n_32893;
wire n_32894;
wire n_32895;
wire n_32896;
wire n_32897;
wire n_32898;
wire n_32899;
wire n_32900;
wire n_32901;
wire n_32902;
wire n_32903;
wire n_32904;
wire n_32905;
wire n_32906;
wire n_32907;
wire n_32908;
wire n_32909;
wire n_32910;
wire n_32911;
wire n_32912;
wire n_32913;
wire n_32914;
wire n_32915;
wire n_32916;
wire n_32917;
wire n_32918;
wire n_32919;
wire n_32920;
wire n_32921;
wire n_32922;
wire n_32923;
wire n_32924;
wire n_32925;
wire n_32926;
wire n_32927;
wire n_32928;
wire n_32929;
wire n_32930;
wire n_32931;
wire n_32932;
wire n_32933;
wire n_32934;
wire n_32935;
wire n_32936;
wire n_32937;
wire n_32938;
wire n_32939;
wire n_32940;
wire n_32941;
wire n_32942;
wire n_32943;
wire n_32944;
wire n_32945;
wire n_32946;
wire n_32947;
wire n_32948;
wire n_32949;
wire n_32950;
wire n_32951;
wire n_32952;
wire n_32953;
wire n_32954;
wire n_32955;
wire n_32956;
wire n_32957;
wire n_32958;
wire n_32959;
wire n_32960;
wire n_32961;
wire n_32962;
wire n_32963;
wire n_32964;
wire n_32965;
wire n_32966;
wire n_32967;
wire n_32968;
wire n_32969;
wire n_32970;
wire n_32971;
wire n_32972;
wire n_32973;
wire n_32974;
wire n_32975;
wire n_32976;
wire n_32977;
wire n_32978;
wire n_32979;
wire n_32980;
wire n_32981;
wire n_32982;
wire n_32983;
wire n_32984;
wire n_32985;
wire n_32986;
wire n_32987;
wire n_32988;
wire n_32989;
wire n_32990;
wire n_32991;
wire n_32992;
wire n_32993;
wire n_32994;
wire n_32995;
wire n_32996;
wire n_32997;
wire n_32998;
wire n_32999;
wire n_33000;
wire n_33001;
wire n_33002;
wire n_33003;
wire n_33004;
wire n_33005;
wire n_33006;
wire n_33007;
wire n_33008;
wire n_33009;
wire n_33010;
wire n_33011;
wire n_33012;
wire n_33013;
wire n_33014;
wire n_33015;
wire n_33016;
wire n_33017;
wire n_33018;
wire n_33019;
wire n_33020;
wire n_33021;
wire n_33022;
wire n_33023;
wire n_33024;
wire n_33025;
wire n_33026;
wire n_33027;
wire n_33028;
wire n_33029;
wire n_33030;
wire n_33031;
wire n_33032;
wire n_33033;
wire n_33034;
wire n_33035;
wire n_33036;
wire n_33037;
wire n_33038;
wire n_33039;
wire n_33040;
wire n_33041;
wire n_33042;
wire n_33043;
wire n_33044;
wire n_33045;
wire n_33046;
wire n_33047;
wire n_33048;
wire n_33049;
wire n_33050;
wire n_33051;
wire n_33052;
wire n_33053;
wire n_33054;
wire n_33055;
wire n_33056;
wire n_33057;
wire n_33058;
wire n_33059;
wire n_33060;
wire n_33061;
wire n_33062;
wire n_33063;
wire n_33064;
wire n_33065;
wire n_33066;
wire n_33067;
wire n_33068;
wire n_33069;
wire n_33070;
wire n_33071;
wire n_33072;
wire n_33073;
wire n_33074;
wire n_33075;
wire n_33076;
wire n_33077;
wire n_33078;
wire n_33079;
wire n_33080;
wire n_33081;
wire n_33082;
wire n_33083;
wire n_33084;
wire n_33085;
wire n_33086;
wire n_33087;
wire n_33088;
wire n_33089;
wire n_33090;
wire n_33091;
wire n_33092;
wire n_33093;
wire n_33094;
wire n_33095;
wire n_33096;
wire n_33097;
wire n_33098;
wire n_33099;
wire n_33100;
wire n_33101;
wire n_33102;
wire n_33103;
wire n_33104;
wire n_33105;
wire n_33106;
wire n_33107;
wire n_33108;
wire n_33109;
wire n_33110;
wire n_33111;
wire n_33112;
wire n_33113;
wire n_33114;
wire n_33115;
wire n_33116;
wire n_33117;
wire n_33118;
wire n_33119;
wire n_33120;
wire n_33121;
wire n_33122;
wire n_33123;
wire n_33124;
wire n_33125;
wire n_33126;
wire n_33127;
wire n_33128;
wire n_33129;
wire n_33130;
wire n_33131;
wire n_33132;
wire n_33133;
wire n_33134;
wire n_33135;
wire n_33136;
wire n_33137;
wire n_33138;
wire n_33139;
wire n_33140;
wire n_33141;
wire n_33142;
wire n_33143;
wire n_33144;
wire n_33145;
wire n_33146;
wire n_33147;
wire n_33148;
wire n_33149;
wire n_33150;
wire n_33151;
wire n_33152;
wire n_33153;
wire n_33154;
wire n_33155;
wire n_33156;
wire n_33157;
wire n_33158;
wire n_33159;
wire n_33160;
wire n_33161;
wire n_33162;
wire n_33163;
wire n_33164;
wire n_33165;
wire n_33166;
wire n_33167;
wire n_33168;
wire n_33169;
wire n_33170;
wire n_33171;
wire n_33172;
wire n_33173;
wire n_33174;
wire n_33175;
wire n_33176;
wire n_33177;
wire n_33178;
wire n_33179;
wire n_33180;
wire n_33181;
wire n_33182;
wire n_33183;
wire n_33184;
wire n_33185;
wire n_33186;
wire n_33187;
wire n_33188;
wire n_33189;
wire n_33190;
wire n_33191;
wire n_33192;
wire n_33193;
wire n_33194;
wire n_33195;
wire n_33196;
wire n_33197;
wire n_33198;
wire n_33199;
wire n_33200;
wire n_33201;
wire n_33202;
wire n_33203;
wire n_33204;
wire n_33205;
wire n_33206;
wire n_33207;
wire n_33208;
wire n_33209;
wire n_33210;
wire n_33211;
wire n_33212;
wire n_33213;
wire n_33214;
wire n_33215;
wire n_33216;
wire n_33217;
wire n_33218;
wire n_33219;
wire n_33220;
wire n_33221;
wire n_33222;
wire n_33223;
wire n_33224;
wire n_33225;
wire n_33226;
wire n_33227;
wire n_33228;
wire n_33229;
wire n_33230;
wire n_33231;
wire n_33232;
wire n_33233;
wire n_33234;
wire n_33235;
wire n_33236;
wire n_33237;
wire n_33238;
wire n_33239;
wire n_33240;
wire n_33241;
wire n_33242;
wire n_33243;
wire n_33244;
wire n_33245;
wire n_33246;
wire n_33247;
wire n_33248;
wire n_33249;
wire n_33250;
wire n_33251;
wire n_33252;
wire n_33253;
wire n_33254;
wire n_33255;
wire n_33256;
wire n_33257;
wire n_33258;
wire n_33259;
wire n_33260;
wire n_33261;
wire n_33262;
wire n_33263;
wire n_33264;
wire n_33265;
wire n_33266;
wire n_33267;
wire n_33268;
wire n_33269;
wire n_33270;
wire n_33271;
wire n_33272;
wire n_33273;
wire n_33274;
wire n_33275;
wire n_33276;
wire n_33277;
wire n_33278;
wire n_33279;
wire n_33280;
wire n_33281;
wire n_33282;
wire n_33283;
wire n_33284;
wire n_33285;
wire n_33286;
wire n_33287;
wire n_33288;
wire n_33289;
wire n_33290;
wire n_33291;
wire n_33292;
wire n_33293;
wire n_33294;
wire n_33295;
wire n_33296;
wire n_33297;
wire n_33298;
wire n_33299;
wire n_33300;
wire n_33301;
wire n_33302;
wire n_33303;
wire n_33304;
wire n_33305;
wire n_33306;
wire n_33307;
wire n_33308;
wire n_33309;
wire n_33310;
wire n_33311;
wire n_33312;
wire n_33313;
wire n_33314;
wire n_33315;
wire n_33316;
wire n_33317;
wire n_33318;
wire n_33319;
wire n_33320;
wire n_33321;
wire n_33322;
wire n_33323;
wire n_33324;
wire n_33325;
wire n_33326;
wire n_33327;
wire n_33328;
wire n_33329;
wire n_33330;
wire n_33331;
wire n_33332;
wire n_33333;
wire n_33334;
wire n_33335;
wire n_33336;
wire n_33337;
wire n_33338;
wire n_33339;
wire n_33340;
wire n_33341;
wire n_33342;
wire n_33343;
wire n_33344;
wire n_33345;
wire n_33346;
wire n_33347;
wire n_33348;
wire n_33349;
wire n_33350;
wire n_33351;
wire n_33352;
wire n_33353;
wire n_33354;
wire n_33355;
wire n_33356;
wire n_33357;
wire n_33358;
wire n_33359;
wire n_33360;
wire n_33361;
wire n_33362;
wire n_33363;
wire n_33364;
wire n_33365;
wire n_33366;
wire n_33367;
wire n_33368;
wire n_33369;
wire n_33370;
wire n_33371;
wire n_33372;
wire n_33373;
wire n_33374;
wire n_33375;
wire n_33376;
wire n_33377;
wire n_33378;
wire n_33379;
wire n_33380;
wire n_33381;
wire n_33382;
wire n_33383;
wire n_33384;
wire n_33385;
wire n_33386;
wire n_33387;
wire n_33388;
wire n_33389;
wire n_33390;
wire n_33391;
wire n_33392;
wire n_33393;
wire n_33394;
wire n_33395;
wire n_33396;
wire n_33397;
wire n_33398;
wire n_33399;
wire n_33400;
wire n_33401;
wire n_33402;
wire n_33403;
wire n_33404;
wire n_33405;
wire n_33406;
wire n_33407;
wire n_33408;
wire n_33409;
wire n_33410;
wire n_33411;
wire n_33412;
wire n_33413;
wire n_33414;
wire n_33415;
wire n_33416;
wire n_33417;
wire n_33418;
wire n_33419;
wire n_33420;
wire n_33421;
wire n_33422;
wire n_33423;
wire n_33424;
wire n_33425;
wire n_33426;
wire n_33427;
wire n_33428;
wire n_33429;
wire n_33430;
wire n_33431;
wire n_33432;
wire n_33433;
wire n_33434;
wire n_33435;
wire n_33436;
wire n_33437;
wire n_33438;
wire n_33439;
wire n_33440;
wire n_33441;
wire n_33442;
wire n_33443;
wire n_33444;
wire n_33445;
wire n_33446;
wire n_33447;
wire n_33448;
wire n_33449;
wire n_33450;
wire n_33451;
wire n_33452;
wire n_33453;
wire n_33454;
wire n_33455;
wire n_33456;
wire n_33457;
wire n_33458;
wire n_33459;
wire n_33460;
wire n_33461;
wire n_33462;
wire n_33463;
wire n_33464;
wire n_33465;
wire n_33466;
wire n_33467;
wire n_33468;
wire n_33469;
wire n_33470;
wire n_33471;
wire n_33472;
wire n_33473;
wire n_33474;
wire n_33475;
wire n_33476;
wire n_33477;
wire n_33478;
wire n_33479;
wire n_33480;
wire n_33481;
wire n_33482;
wire n_33483;
wire n_33484;
wire n_33485;
wire n_33486;
wire n_33487;
wire n_33488;
wire n_33489;
wire n_33490;
wire n_33491;
wire n_33492;
wire n_33493;
wire n_33494;
wire n_33495;
wire n_33496;
wire n_33497;
wire n_33498;
wire n_33499;
wire n_33500;
wire n_33501;
wire n_33502;
wire n_33503;
wire n_33504;
wire n_33505;
wire n_33506;
wire n_33507;
wire n_33508;
wire n_33509;
wire n_33510;
wire n_33511;
wire n_33512;
wire n_33513;
wire n_33514;
wire n_33515;
wire n_33516;
wire n_33517;
wire n_33518;
wire n_33519;
wire n_33520;
wire n_33521;
wire n_33522;
wire n_33523;
wire n_33524;
wire n_33525;
wire n_33526;
wire n_33527;
wire n_33528;
wire n_33529;
wire n_33530;
wire n_33531;
wire n_33532;
wire n_33533;
wire n_33534;
wire n_33535;
wire n_33536;
wire n_33537;
wire n_33538;
wire n_33539;
wire n_33540;
wire n_33541;
wire n_33542;
wire n_33543;
wire n_33544;
wire n_33545;
wire n_33546;
wire n_33547;
wire n_33548;
wire n_33549;
wire n_33550;
wire n_33551;
wire n_33552;
wire n_33553;
wire n_33554;
wire n_33555;
wire n_33556;
wire n_33557;
wire n_33558;
wire n_33559;
wire n_33560;
wire n_33561;
wire n_33562;
wire n_33563;
wire n_33564;
wire n_33565;
wire n_33566;
wire n_33567;
wire n_33568;
wire n_33569;
wire n_33570;
wire n_33571;
wire n_33572;
wire n_33573;
wire n_33574;
wire n_33575;
wire n_33576;
wire n_33577;
wire n_33578;
wire n_33579;
wire n_33580;
wire n_33581;
wire n_33582;
wire n_33583;
wire n_33584;
wire n_33585;
wire n_33586;
wire n_33587;
wire n_33588;
wire n_33589;
wire n_33590;
wire n_33591;
wire n_33592;
wire n_33593;
wire n_33594;
wire n_33595;
wire n_33596;
wire n_33597;
wire n_33598;
wire n_33599;
wire n_33600;
wire n_33601;
wire n_33602;
wire n_33603;
wire n_33604;
wire n_33605;
wire n_33606;
wire n_33607;
wire n_33608;
wire n_33609;
wire n_33610;
wire n_33611;
wire n_33612;
wire n_33613;
wire n_33614;
wire n_33615;
wire n_33616;
wire n_33617;
wire n_33618;
wire n_33619;
wire n_33620;
wire n_33621;
wire n_33622;
wire n_33623;
wire n_33624;
wire n_33625;
wire n_33626;
wire n_33627;
wire n_33628;
wire n_33629;
wire n_33630;
wire n_33631;
wire n_33632;
wire n_33633;
wire n_33634;
wire n_33635;
wire n_33636;
wire n_33637;
wire n_33638;
wire n_33639;
wire n_33640;
wire n_33641;
wire n_33642;
wire n_33643;
wire n_33644;
wire n_33645;
wire n_33646;
wire n_33647;
wire n_33648;
wire n_33649;
wire n_33650;
wire n_33651;
wire n_33652;
wire n_33653;
wire n_33654;
wire n_33655;
wire n_33656;
wire n_33657;
wire n_33658;
wire n_33659;
wire n_33660;
wire n_33661;
wire n_33662;
wire n_33663;
wire n_33664;
wire n_33665;
wire n_33666;
wire n_33667;
wire n_33668;
wire n_33669;
wire n_33670;
wire n_33671;
wire n_33672;
wire n_33673;
wire n_33674;
wire n_33675;
wire n_33676;
wire n_33677;
wire n_33678;
wire n_33679;
wire n_33680;
wire n_33681;
wire n_33682;
wire n_33683;
wire n_33684;
wire n_33685;
wire n_33686;
wire n_33687;
wire n_33688;
wire n_33689;
wire n_33690;
wire n_33691;
wire n_33692;
wire n_33693;
wire n_33694;
wire n_33695;
wire n_33696;
wire n_33697;
wire n_33698;
wire n_33699;
wire n_33700;
wire n_33701;
wire n_33702;
wire n_33703;
wire n_33704;
wire n_33705;
wire n_33706;
wire n_33707;
wire n_33708;
wire n_33709;
wire n_33710;
wire n_33711;
wire n_33712;
wire n_33713;
wire n_33714;
wire n_33715;
wire n_33716;
wire n_33717;
wire n_33718;
wire n_33719;
wire n_33720;
wire n_33721;
wire n_33722;
wire n_33723;
wire n_33724;
wire n_33725;
wire n_33726;
wire n_33727;
wire n_33728;
wire n_33729;
wire n_33730;
wire n_33731;
wire n_33732;
wire n_33733;
wire n_33734;
wire n_33735;
wire n_33736;
wire n_33737;
wire n_33738;
wire n_33739;
wire n_33740;
wire n_33741;
wire n_33742;
wire n_33743;
wire n_33744;
wire n_33745;
wire n_33746;
wire n_33747;
wire n_33748;
wire n_33749;
wire n_33750;
wire n_33751;
wire n_33752;
wire n_33753;
wire n_33754;
wire n_33755;
wire n_33756;
wire n_33757;
wire n_33758;
wire n_33759;
wire n_33760;
wire n_33761;
wire n_33762;
wire n_33763;
wire n_33764;
wire n_33765;
wire n_33766;
wire n_33767;
wire n_33768;
wire n_33769;
wire n_33770;
wire n_33771;
wire n_33772;
wire n_33773;
wire n_33774;
wire n_33775;
wire n_33776;
wire n_33777;
wire n_33778;
wire n_33779;
wire n_33780;
wire n_33781;
wire n_33782;
wire n_33783;
wire n_33784;
wire n_33785;
wire n_33786;
wire n_33787;
wire n_33788;
wire n_33789;
wire n_33790;
wire n_33791;
wire n_33792;
wire n_33793;
wire n_33794;
wire n_33795;
wire n_33796;
wire n_33797;
wire n_33798;
wire n_33799;
wire n_33800;
wire n_33801;
wire n_33802;
wire n_33803;
wire n_33804;
wire n_33805;
wire n_33806;
wire n_33807;
wire n_33808;
wire n_33809;
wire n_33810;
wire n_33811;
wire n_33812;
wire n_33813;
wire n_33814;
wire n_33815;
wire n_33816;
wire n_33817;
wire n_33818;
wire n_33819;
wire n_33820;
wire n_33821;
wire n_33822;
wire n_33823;
wire n_33824;
wire n_33825;
assign n_1 = ~x_40 &  x_41;
assign n_2 =  x_42 &  n_1;
assign n_3 =  x_39 &  n_2;
assign n_4 = ~x_37 &  x_38;
assign n_5 = ~x_33 &  x_34;
assign n_6 =  x_35 &  n_5;
assign n_7 = ~x_36 &  n_6;
assign n_8 =  n_4 &  n_7;
assign n_9 =  n_3 &  n_8;
assign n_10 =  x_2375 & ~n_9;
assign n_11 =  i_29 &  n_9;
assign n_12 = ~n_10 & ~n_11;
assign n_13 =  x_2375 & ~n_12;
assign n_14 = ~x_2375 &  n_12;
assign n_15 = ~n_13 & ~n_14;
assign n_16 =  x_2374 & ~n_9;
assign n_17 =  i_28 &  n_9;
assign n_18 = ~n_16 & ~n_17;
assign n_19 =  x_2374 & ~n_18;
assign n_20 = ~x_2374 &  n_18;
assign n_21 = ~n_19 & ~n_20;
assign n_22 =  x_2373 & ~n_9;
assign n_23 =  i_27 &  n_9;
assign n_24 = ~n_22 & ~n_23;
assign n_25 =  x_2373 & ~n_24;
assign n_26 = ~x_2373 &  n_24;
assign n_27 = ~n_25 & ~n_26;
assign n_28 =  x_2372 & ~n_9;
assign n_29 =  i_26 &  n_9;
assign n_30 = ~n_28 & ~n_29;
assign n_31 =  x_2372 & ~n_30;
assign n_32 = ~x_2372 &  n_30;
assign n_33 = ~n_31 & ~n_32;
assign n_34 =  x_2371 & ~n_9;
assign n_35 =  i_25 &  n_9;
assign n_36 = ~n_34 & ~n_35;
assign n_37 =  x_2371 & ~n_36;
assign n_38 = ~x_2371 &  n_36;
assign n_39 = ~n_37 & ~n_38;
assign n_40 =  x_2370 & ~n_9;
assign n_41 =  i_24 &  n_9;
assign n_42 = ~n_40 & ~n_41;
assign n_43 =  x_2370 & ~n_42;
assign n_44 = ~x_2370 &  n_42;
assign n_45 = ~n_43 & ~n_44;
assign n_46 =  x_2369 & ~n_9;
assign n_47 =  i_23 &  n_9;
assign n_48 = ~n_46 & ~n_47;
assign n_49 =  x_2369 & ~n_48;
assign n_50 = ~x_2369 &  n_48;
assign n_51 = ~n_49 & ~n_50;
assign n_52 =  x_2368 & ~n_9;
assign n_53 =  i_22 &  n_9;
assign n_54 = ~n_52 & ~n_53;
assign n_55 =  x_2368 & ~n_54;
assign n_56 = ~x_2368 &  n_54;
assign n_57 = ~n_55 & ~n_56;
assign n_58 =  x_2367 & ~n_9;
assign n_59 =  i_21 &  n_9;
assign n_60 = ~n_58 & ~n_59;
assign n_61 =  x_2367 & ~n_60;
assign n_62 = ~x_2367 &  n_60;
assign n_63 = ~n_61 & ~n_62;
assign n_64 =  x_2366 & ~n_9;
assign n_65 =  i_20 &  n_9;
assign n_66 = ~n_64 & ~n_65;
assign n_67 =  x_2366 & ~n_66;
assign n_68 = ~x_2366 &  n_66;
assign n_69 = ~n_67 & ~n_68;
assign n_70 =  x_2365 & ~n_9;
assign n_71 =  i_19 &  n_9;
assign n_72 = ~n_70 & ~n_71;
assign n_73 =  x_2365 & ~n_72;
assign n_74 = ~x_2365 &  n_72;
assign n_75 = ~n_73 & ~n_74;
assign n_76 =  x_2364 & ~n_9;
assign n_77 =  i_18 &  n_9;
assign n_78 = ~n_76 & ~n_77;
assign n_79 =  x_2364 & ~n_78;
assign n_80 = ~x_2364 &  n_78;
assign n_81 = ~n_79 & ~n_80;
assign n_82 =  x_2363 & ~n_9;
assign n_83 =  i_17 &  n_9;
assign n_84 = ~n_82 & ~n_83;
assign n_85 =  x_2363 & ~n_84;
assign n_86 = ~x_2363 &  n_84;
assign n_87 = ~n_85 & ~n_86;
assign n_88 =  x_2362 & ~n_9;
assign n_89 =  i_16 &  n_9;
assign n_90 = ~n_88 & ~n_89;
assign n_91 =  x_2362 & ~n_90;
assign n_92 = ~x_2362 &  n_90;
assign n_93 = ~n_91 & ~n_92;
assign n_94 =  x_2361 & ~n_9;
assign n_95 =  i_15 &  n_9;
assign n_96 = ~n_94 & ~n_95;
assign n_97 =  x_2361 & ~n_96;
assign n_98 = ~x_2361 &  n_96;
assign n_99 = ~n_97 & ~n_98;
assign n_100 =  x_2360 & ~n_9;
assign n_101 =  i_14 &  n_9;
assign n_102 = ~n_100 & ~n_101;
assign n_103 =  x_2360 & ~n_102;
assign n_104 = ~x_2360 &  n_102;
assign n_105 = ~n_103 & ~n_104;
assign n_106 =  x_2359 & ~n_9;
assign n_107 =  i_13 &  n_9;
assign n_108 = ~n_106 & ~n_107;
assign n_109 =  x_2359 & ~n_108;
assign n_110 = ~x_2359 &  n_108;
assign n_111 = ~n_109 & ~n_110;
assign n_112 =  x_2358 & ~n_9;
assign n_113 =  i_12 &  n_9;
assign n_114 = ~n_112 & ~n_113;
assign n_115 =  x_2358 & ~n_114;
assign n_116 = ~x_2358 &  n_114;
assign n_117 = ~n_115 & ~n_116;
assign n_118 =  x_2357 & ~n_9;
assign n_119 =  i_11 &  n_9;
assign n_120 = ~n_118 & ~n_119;
assign n_121 =  x_2357 & ~n_120;
assign n_122 = ~x_2357 &  n_120;
assign n_123 = ~n_121 & ~n_122;
assign n_124 =  x_2356 & ~n_9;
assign n_125 =  i_10 &  n_9;
assign n_126 = ~n_124 & ~n_125;
assign n_127 =  x_2356 & ~n_126;
assign n_128 = ~x_2356 &  n_126;
assign n_129 = ~n_127 & ~n_128;
assign n_130 =  x_2355 & ~n_9;
assign n_131 =  i_9 &  n_9;
assign n_132 = ~n_130 & ~n_131;
assign n_133 =  x_2355 & ~n_132;
assign n_134 = ~x_2355 &  n_132;
assign n_135 = ~n_133 & ~n_134;
assign n_136 =  x_2354 & ~n_9;
assign n_137 =  i_8 &  n_9;
assign n_138 = ~n_136 & ~n_137;
assign n_139 =  x_2354 & ~n_138;
assign n_140 = ~x_2354 &  n_138;
assign n_141 = ~n_139 & ~n_140;
assign n_142 =  x_2353 & ~n_9;
assign n_143 =  i_7 &  n_9;
assign n_144 = ~n_142 & ~n_143;
assign n_145 =  x_2353 & ~n_144;
assign n_146 = ~x_2353 &  n_144;
assign n_147 = ~n_145 & ~n_146;
assign n_148 =  x_2352 & ~n_9;
assign n_149 =  i_6 &  n_9;
assign n_150 = ~n_148 & ~n_149;
assign n_151 =  x_2352 & ~n_150;
assign n_152 = ~x_2352 &  n_150;
assign n_153 = ~n_151 & ~n_152;
assign n_154 =  x_2351 & ~n_9;
assign n_155 =  i_5 &  n_9;
assign n_156 = ~n_154 & ~n_155;
assign n_157 =  x_2351 & ~n_156;
assign n_158 = ~x_2351 &  n_156;
assign n_159 = ~n_157 & ~n_158;
assign n_160 =  x_2350 & ~n_9;
assign n_161 =  i_4 &  n_9;
assign n_162 = ~n_160 & ~n_161;
assign n_163 =  x_2350 & ~n_162;
assign n_164 = ~x_2350 &  n_162;
assign n_165 = ~n_163 & ~n_164;
assign n_166 =  x_2349 & ~n_9;
assign n_167 =  i_3 &  n_9;
assign n_168 = ~n_166 & ~n_167;
assign n_169 =  x_2349 & ~n_168;
assign n_170 = ~x_2349 &  n_168;
assign n_171 = ~n_169 & ~n_170;
assign n_172 =  x_2348 & ~n_9;
assign n_173 =  i_2 &  n_9;
assign n_174 = ~n_172 & ~n_173;
assign n_175 =  x_2348 & ~n_174;
assign n_176 = ~x_2348 &  n_174;
assign n_177 = ~n_175 & ~n_176;
assign n_178 =  x_2347 & ~n_9;
assign n_179 =  i_1 &  n_9;
assign n_180 = ~n_178 & ~n_179;
assign n_181 =  x_2347 & ~n_180;
assign n_182 = ~x_2347 &  n_180;
assign n_183 = ~n_181 & ~n_182;
assign n_184 = ~x_39 & ~x_40;
assign n_185 =  x_41 & ~x_42;
assign n_186 =  n_184 &  n_185;
assign n_187 =  x_37 & ~x_38;
assign n_188 = ~x_35 &  x_36;
assign n_189 = ~x_33 & ~x_34;
assign n_190 =  n_188 &  n_189;
assign n_191 =  n_187 &  n_190;
assign n_192 =  n_186 &  n_191;
assign n_193 =  x_2346 & ~n_192;
assign n_194 =  i_32 &  n_192;
assign n_195 = ~n_193 & ~n_194;
assign n_196 =  x_2346 & ~n_195;
assign n_197 = ~x_2346 &  n_195;
assign n_198 = ~n_196 & ~n_197;
assign n_199 =  x_2345 & ~n_192;
assign n_200 =  i_31 &  n_192;
assign n_201 = ~n_199 & ~n_200;
assign n_202 =  x_2345 & ~n_201;
assign n_203 = ~x_2345 &  n_201;
assign n_204 = ~n_202 & ~n_203;
assign n_205 =  x_2344 & ~n_192;
assign n_206 =  i_30 &  n_192;
assign n_207 = ~n_205 & ~n_206;
assign n_208 =  x_2344 & ~n_207;
assign n_209 = ~x_2344 &  n_207;
assign n_210 = ~n_208 & ~n_209;
assign n_211 =  x_2343 & ~n_192;
assign n_212 =  i_29 &  n_192;
assign n_213 = ~n_211 & ~n_212;
assign n_214 =  x_2343 & ~n_213;
assign n_215 = ~x_2343 &  n_213;
assign n_216 = ~n_214 & ~n_215;
assign n_217 =  x_2342 & ~n_192;
assign n_218 =  i_28 &  n_192;
assign n_219 = ~n_217 & ~n_218;
assign n_220 =  x_2342 & ~n_219;
assign n_221 = ~x_2342 &  n_219;
assign n_222 = ~n_220 & ~n_221;
assign n_223 =  x_2341 & ~n_192;
assign n_224 =  i_27 &  n_192;
assign n_225 = ~n_223 & ~n_224;
assign n_226 =  x_2341 & ~n_225;
assign n_227 = ~x_2341 &  n_225;
assign n_228 = ~n_226 & ~n_227;
assign n_229 =  x_2340 & ~n_192;
assign n_230 =  i_26 &  n_192;
assign n_231 = ~n_229 & ~n_230;
assign n_232 =  x_2340 & ~n_231;
assign n_233 = ~x_2340 &  n_231;
assign n_234 = ~n_232 & ~n_233;
assign n_235 =  x_2339 & ~n_192;
assign n_236 =  i_25 &  n_192;
assign n_237 = ~n_235 & ~n_236;
assign n_238 =  x_2339 & ~n_237;
assign n_239 = ~x_2339 &  n_237;
assign n_240 = ~n_238 & ~n_239;
assign n_241 =  x_2338 & ~n_192;
assign n_242 =  i_24 &  n_192;
assign n_243 = ~n_241 & ~n_242;
assign n_244 =  x_2338 & ~n_243;
assign n_245 = ~x_2338 &  n_243;
assign n_246 = ~n_244 & ~n_245;
assign n_247 =  x_2337 & ~n_192;
assign n_248 =  i_23 &  n_192;
assign n_249 = ~n_247 & ~n_248;
assign n_250 =  x_2337 & ~n_249;
assign n_251 = ~x_2337 &  n_249;
assign n_252 = ~n_250 & ~n_251;
assign n_253 =  x_2336 & ~n_192;
assign n_254 =  i_22 &  n_192;
assign n_255 = ~n_253 & ~n_254;
assign n_256 =  x_2336 & ~n_255;
assign n_257 = ~x_2336 &  n_255;
assign n_258 = ~n_256 & ~n_257;
assign n_259 =  x_2335 & ~n_192;
assign n_260 =  i_21 &  n_192;
assign n_261 = ~n_259 & ~n_260;
assign n_262 =  x_2335 & ~n_261;
assign n_263 = ~x_2335 &  n_261;
assign n_264 = ~n_262 & ~n_263;
assign n_265 =  x_2334 & ~n_192;
assign n_266 =  i_20 &  n_192;
assign n_267 = ~n_265 & ~n_266;
assign n_268 =  x_2334 & ~n_267;
assign n_269 = ~x_2334 &  n_267;
assign n_270 = ~n_268 & ~n_269;
assign n_271 =  x_2333 & ~n_192;
assign n_272 =  i_19 &  n_192;
assign n_273 = ~n_271 & ~n_272;
assign n_274 =  x_2333 & ~n_273;
assign n_275 = ~x_2333 &  n_273;
assign n_276 = ~n_274 & ~n_275;
assign n_277 =  x_2332 & ~n_192;
assign n_278 =  i_18 &  n_192;
assign n_279 = ~n_277 & ~n_278;
assign n_280 =  x_2332 & ~n_279;
assign n_281 = ~x_2332 &  n_279;
assign n_282 = ~n_280 & ~n_281;
assign n_283 =  x_2331 & ~n_192;
assign n_284 =  i_17 &  n_192;
assign n_285 = ~n_283 & ~n_284;
assign n_286 =  x_2331 & ~n_285;
assign n_287 = ~x_2331 &  n_285;
assign n_288 = ~n_286 & ~n_287;
assign n_289 =  x_2330 & ~n_192;
assign n_290 =  i_16 &  n_192;
assign n_291 = ~n_289 & ~n_290;
assign n_292 =  x_2330 & ~n_291;
assign n_293 = ~x_2330 &  n_291;
assign n_294 = ~n_292 & ~n_293;
assign n_295 =  x_2329 & ~n_192;
assign n_296 =  i_15 &  n_192;
assign n_297 = ~n_295 & ~n_296;
assign n_298 =  x_2329 & ~n_297;
assign n_299 = ~x_2329 &  n_297;
assign n_300 = ~n_298 & ~n_299;
assign n_301 =  x_2328 & ~n_192;
assign n_302 =  i_14 &  n_192;
assign n_303 = ~n_301 & ~n_302;
assign n_304 =  x_2328 & ~n_303;
assign n_305 = ~x_2328 &  n_303;
assign n_306 = ~n_304 & ~n_305;
assign n_307 =  x_2327 & ~n_192;
assign n_308 =  i_13 &  n_192;
assign n_309 = ~n_307 & ~n_308;
assign n_310 =  x_2327 & ~n_309;
assign n_311 = ~x_2327 &  n_309;
assign n_312 = ~n_310 & ~n_311;
assign n_313 =  x_2326 & ~n_192;
assign n_314 =  i_12 &  n_192;
assign n_315 = ~n_313 & ~n_314;
assign n_316 =  x_2326 & ~n_315;
assign n_317 = ~x_2326 &  n_315;
assign n_318 = ~n_316 & ~n_317;
assign n_319 =  x_2325 & ~n_192;
assign n_320 =  i_11 &  n_192;
assign n_321 = ~n_319 & ~n_320;
assign n_322 =  x_2325 & ~n_321;
assign n_323 = ~x_2325 &  n_321;
assign n_324 = ~n_322 & ~n_323;
assign n_325 =  x_2324 & ~n_192;
assign n_326 =  i_10 &  n_192;
assign n_327 = ~n_325 & ~n_326;
assign n_328 =  x_2324 & ~n_327;
assign n_329 = ~x_2324 &  n_327;
assign n_330 = ~n_328 & ~n_329;
assign n_331 =  x_2323 & ~n_192;
assign n_332 =  i_9 &  n_192;
assign n_333 = ~n_331 & ~n_332;
assign n_334 =  x_2323 & ~n_333;
assign n_335 = ~x_2323 &  n_333;
assign n_336 = ~n_334 & ~n_335;
assign n_337 =  x_2322 & ~n_192;
assign n_338 =  i_8 &  n_192;
assign n_339 = ~n_337 & ~n_338;
assign n_340 =  x_2322 & ~n_339;
assign n_341 = ~x_2322 &  n_339;
assign n_342 = ~n_340 & ~n_341;
assign n_343 =  x_2321 & ~n_192;
assign n_344 =  i_7 &  n_192;
assign n_345 = ~n_343 & ~n_344;
assign n_346 =  x_2321 & ~n_345;
assign n_347 = ~x_2321 &  n_345;
assign n_348 = ~n_346 & ~n_347;
assign n_349 =  x_2320 & ~n_192;
assign n_350 =  i_6 &  n_192;
assign n_351 = ~n_349 & ~n_350;
assign n_352 =  x_2320 & ~n_351;
assign n_353 = ~x_2320 &  n_351;
assign n_354 = ~n_352 & ~n_353;
assign n_355 =  x_2319 & ~n_192;
assign n_356 =  i_5 &  n_192;
assign n_357 = ~n_355 & ~n_356;
assign n_358 =  x_2319 & ~n_357;
assign n_359 = ~x_2319 &  n_357;
assign n_360 = ~n_358 & ~n_359;
assign n_361 =  x_2318 & ~n_192;
assign n_362 =  i_4 &  n_192;
assign n_363 = ~n_361 & ~n_362;
assign n_364 =  x_2318 & ~n_363;
assign n_365 = ~x_2318 &  n_363;
assign n_366 = ~n_364 & ~n_365;
assign n_367 =  x_2317 & ~n_192;
assign n_368 =  i_3 &  n_192;
assign n_369 = ~n_367 & ~n_368;
assign n_370 =  x_2317 & ~n_369;
assign n_371 = ~x_2317 &  n_369;
assign n_372 = ~n_370 & ~n_371;
assign n_373 =  x_2316 & ~n_192;
assign n_374 =  i_2 &  n_192;
assign n_375 = ~n_373 & ~n_374;
assign n_376 =  x_2316 & ~n_375;
assign n_377 = ~x_2316 &  n_375;
assign n_378 = ~n_376 & ~n_377;
assign n_379 =  x_2315 & ~n_192;
assign n_380 =  i_1 &  n_192;
assign n_381 = ~n_379 & ~n_380;
assign n_382 =  x_2315 & ~n_381;
assign n_383 = ~x_2315 &  n_381;
assign n_384 = ~n_382 & ~n_383;
assign n_385 =  x_39 & ~x_40;
assign n_386 = ~x_42 &  n_385;
assign n_387 = ~x_35 &  n_5;
assign n_388 =  x_36 &  n_387;
assign n_389 =  x_37 &  x_38;
assign n_390 =  n_388 &  n_389;
assign n_391 =  n_386 &  n_390;
assign n_392 = ~x_41 &  n_391;
assign n_393 =  x_2314 & ~n_392;
assign n_394 =  i_32 &  n_392;
assign n_395 = ~n_393 & ~n_394;
assign n_396 =  x_2314 & ~n_395;
assign n_397 = ~x_2314 &  n_395;
assign n_398 = ~n_396 & ~n_397;
assign n_399 =  x_2313 & ~n_392;
assign n_400 =  i_31 &  n_392;
assign n_401 = ~n_399 & ~n_400;
assign n_402 =  x_2313 & ~n_401;
assign n_403 = ~x_2313 &  n_401;
assign n_404 = ~n_402 & ~n_403;
assign n_405 =  x_2312 & ~n_392;
assign n_406 =  i_30 &  n_392;
assign n_407 = ~n_405 & ~n_406;
assign n_408 =  x_2312 & ~n_407;
assign n_409 = ~x_2312 &  n_407;
assign n_410 = ~n_408 & ~n_409;
assign n_411 =  x_2311 & ~n_392;
assign n_412 =  i_29 &  n_392;
assign n_413 = ~n_411 & ~n_412;
assign n_414 =  x_2311 & ~n_413;
assign n_415 = ~x_2311 &  n_413;
assign n_416 = ~n_414 & ~n_415;
assign n_417 =  x_2310 & ~n_392;
assign n_418 =  i_28 &  n_392;
assign n_419 = ~n_417 & ~n_418;
assign n_420 =  x_2310 & ~n_419;
assign n_421 = ~x_2310 &  n_419;
assign n_422 = ~n_420 & ~n_421;
assign n_423 =  x_2309 & ~n_392;
assign n_424 =  i_27 &  n_392;
assign n_425 = ~n_423 & ~n_424;
assign n_426 =  x_2309 & ~n_425;
assign n_427 = ~x_2309 &  n_425;
assign n_428 = ~n_426 & ~n_427;
assign n_429 =  x_2308 & ~n_392;
assign n_430 =  i_26 &  n_392;
assign n_431 = ~n_429 & ~n_430;
assign n_432 =  x_2308 & ~n_431;
assign n_433 = ~x_2308 &  n_431;
assign n_434 = ~n_432 & ~n_433;
assign n_435 =  x_2307 & ~n_392;
assign n_436 =  i_25 &  n_392;
assign n_437 = ~n_435 & ~n_436;
assign n_438 =  x_2307 & ~n_437;
assign n_439 = ~x_2307 &  n_437;
assign n_440 = ~n_438 & ~n_439;
assign n_441 =  x_2306 & ~n_392;
assign n_442 =  i_24 &  n_392;
assign n_443 = ~n_441 & ~n_442;
assign n_444 =  x_2306 & ~n_443;
assign n_445 = ~x_2306 &  n_443;
assign n_446 = ~n_444 & ~n_445;
assign n_447 =  x_2305 & ~n_392;
assign n_448 =  i_23 &  n_392;
assign n_449 = ~n_447 & ~n_448;
assign n_450 =  x_2305 & ~n_449;
assign n_451 = ~x_2305 &  n_449;
assign n_452 = ~n_450 & ~n_451;
assign n_453 =  x_2304 & ~n_392;
assign n_454 =  i_22 &  n_392;
assign n_455 = ~n_453 & ~n_454;
assign n_456 =  x_2304 & ~n_455;
assign n_457 = ~x_2304 &  n_455;
assign n_458 = ~n_456 & ~n_457;
assign n_459 =  x_2303 & ~n_392;
assign n_460 =  i_21 &  n_392;
assign n_461 = ~n_459 & ~n_460;
assign n_462 =  x_2303 & ~n_461;
assign n_463 = ~x_2303 &  n_461;
assign n_464 = ~n_462 & ~n_463;
assign n_465 =  x_2302 & ~n_392;
assign n_466 =  i_20 &  n_392;
assign n_467 = ~n_465 & ~n_466;
assign n_468 =  x_2302 & ~n_467;
assign n_469 = ~x_2302 &  n_467;
assign n_470 = ~n_468 & ~n_469;
assign n_471 =  x_2301 & ~n_392;
assign n_472 =  i_19 &  n_392;
assign n_473 = ~n_471 & ~n_472;
assign n_474 =  x_2301 & ~n_473;
assign n_475 = ~x_2301 &  n_473;
assign n_476 = ~n_474 & ~n_475;
assign n_477 =  x_2300 & ~n_392;
assign n_478 =  i_18 &  n_392;
assign n_479 = ~n_477 & ~n_478;
assign n_480 =  x_2300 & ~n_479;
assign n_481 = ~x_2300 &  n_479;
assign n_482 = ~n_480 & ~n_481;
assign n_483 =  x_2299 & ~n_392;
assign n_484 =  i_17 &  n_392;
assign n_485 = ~n_483 & ~n_484;
assign n_486 =  x_2299 & ~n_485;
assign n_487 = ~x_2299 &  n_485;
assign n_488 = ~n_486 & ~n_487;
assign n_489 =  x_2298 & ~n_392;
assign n_490 =  i_16 &  n_392;
assign n_491 = ~n_489 & ~n_490;
assign n_492 =  x_2298 & ~n_491;
assign n_493 = ~x_2298 &  n_491;
assign n_494 = ~n_492 & ~n_493;
assign n_495 =  x_2297 & ~n_392;
assign n_496 =  i_15 &  n_392;
assign n_497 = ~n_495 & ~n_496;
assign n_498 =  x_2297 & ~n_497;
assign n_499 = ~x_2297 &  n_497;
assign n_500 = ~n_498 & ~n_499;
assign n_501 =  x_2296 & ~n_392;
assign n_502 =  i_14 &  n_392;
assign n_503 = ~n_501 & ~n_502;
assign n_504 =  x_2296 & ~n_503;
assign n_505 = ~x_2296 &  n_503;
assign n_506 = ~n_504 & ~n_505;
assign n_507 =  x_2295 & ~n_392;
assign n_508 =  i_13 &  n_392;
assign n_509 = ~n_507 & ~n_508;
assign n_510 =  x_2295 & ~n_509;
assign n_511 = ~x_2295 &  n_509;
assign n_512 = ~n_510 & ~n_511;
assign n_513 =  x_2294 & ~n_392;
assign n_514 =  i_12 &  n_392;
assign n_515 = ~n_513 & ~n_514;
assign n_516 =  x_2294 & ~n_515;
assign n_517 = ~x_2294 &  n_515;
assign n_518 = ~n_516 & ~n_517;
assign n_519 =  x_2293 & ~n_392;
assign n_520 =  i_11 &  n_392;
assign n_521 = ~n_519 & ~n_520;
assign n_522 =  x_2293 & ~n_521;
assign n_523 = ~x_2293 &  n_521;
assign n_524 = ~n_522 & ~n_523;
assign n_525 =  x_2292 & ~n_392;
assign n_526 =  i_10 &  n_392;
assign n_527 = ~n_525 & ~n_526;
assign n_528 =  x_2292 & ~n_527;
assign n_529 = ~x_2292 &  n_527;
assign n_530 = ~n_528 & ~n_529;
assign n_531 =  x_2291 & ~n_392;
assign n_532 =  i_9 &  n_392;
assign n_533 = ~n_531 & ~n_532;
assign n_534 =  x_2291 & ~n_533;
assign n_535 = ~x_2291 &  n_533;
assign n_536 = ~n_534 & ~n_535;
assign n_537 =  x_2290 & ~n_392;
assign n_538 =  i_8 &  n_392;
assign n_539 = ~n_537 & ~n_538;
assign n_540 =  x_2290 & ~n_539;
assign n_541 = ~x_2290 &  n_539;
assign n_542 = ~n_540 & ~n_541;
assign n_543 =  x_2289 & ~n_392;
assign n_544 =  i_7 &  n_392;
assign n_545 = ~n_543 & ~n_544;
assign n_546 =  x_2289 & ~n_545;
assign n_547 = ~x_2289 &  n_545;
assign n_548 = ~n_546 & ~n_547;
assign n_549 =  x_2288 & ~n_392;
assign n_550 =  i_6 &  n_392;
assign n_551 = ~n_549 & ~n_550;
assign n_552 =  x_2288 & ~n_551;
assign n_553 = ~x_2288 &  n_551;
assign n_554 = ~n_552 & ~n_553;
assign n_555 =  x_2287 & ~n_392;
assign n_556 =  i_5 &  n_392;
assign n_557 = ~n_555 & ~n_556;
assign n_558 =  x_2287 & ~n_557;
assign n_559 = ~x_2287 &  n_557;
assign n_560 = ~n_558 & ~n_559;
assign n_561 =  x_2286 & ~n_392;
assign n_562 =  i_4 &  n_392;
assign n_563 = ~n_561 & ~n_562;
assign n_564 =  x_2286 & ~n_563;
assign n_565 = ~x_2286 &  n_563;
assign n_566 = ~n_564 & ~n_565;
assign n_567 =  x_2285 & ~n_392;
assign n_568 =  i_3 &  n_392;
assign n_569 = ~n_567 & ~n_568;
assign n_570 =  x_2285 & ~n_569;
assign n_571 = ~x_2285 &  n_569;
assign n_572 = ~n_570 & ~n_571;
assign n_573 =  x_2284 & ~n_392;
assign n_574 =  i_2 &  n_392;
assign n_575 = ~n_573 & ~n_574;
assign n_576 =  x_2284 & ~n_575;
assign n_577 = ~x_2284 &  n_575;
assign n_578 = ~n_576 & ~n_577;
assign n_579 =  x_2283 & ~n_392;
assign n_580 =  i_1 &  n_392;
assign n_581 = ~n_579 & ~n_580;
assign n_582 =  x_2283 & ~n_581;
assign n_583 = ~x_2283 &  n_581;
assign n_584 = ~n_582 & ~n_583;
assign n_585 =  x_40 & ~x_41;
assign n_586 =  x_42 &  n_585;
assign n_587 =  x_39 &  n_586;
assign n_588 =  n_388 &  n_4;
assign n_589 =  n_587 &  n_588;
assign n_590 =  x_2282 & ~n_589;
assign n_591 =  i_32 &  n_589;
assign n_592 = ~n_590 & ~n_591;
assign n_593 =  x_2282 & ~n_592;
assign n_594 = ~x_2282 &  n_592;
assign n_595 = ~n_593 & ~n_594;
assign n_596 =  x_2281 & ~n_589;
assign n_597 =  i_31 &  n_589;
assign n_598 = ~n_596 & ~n_597;
assign n_599 =  x_2281 & ~n_598;
assign n_600 = ~x_2281 &  n_598;
assign n_601 = ~n_599 & ~n_600;
assign n_602 =  x_2280 & ~n_589;
assign n_603 =  i_30 &  n_589;
assign n_604 = ~n_602 & ~n_603;
assign n_605 =  x_2280 & ~n_604;
assign n_606 = ~x_2280 &  n_604;
assign n_607 = ~n_605 & ~n_606;
assign n_608 =  x_2279 & ~n_589;
assign n_609 =  i_29 &  n_589;
assign n_610 = ~n_608 & ~n_609;
assign n_611 =  x_2279 & ~n_610;
assign n_612 = ~x_2279 &  n_610;
assign n_613 = ~n_611 & ~n_612;
assign n_614 =  x_2278 & ~n_589;
assign n_615 =  i_28 &  n_589;
assign n_616 = ~n_614 & ~n_615;
assign n_617 =  x_2278 & ~n_616;
assign n_618 = ~x_2278 &  n_616;
assign n_619 = ~n_617 & ~n_618;
assign n_620 =  x_2277 & ~n_589;
assign n_621 =  i_27 &  n_589;
assign n_622 = ~n_620 & ~n_621;
assign n_623 =  x_2277 & ~n_622;
assign n_624 = ~x_2277 &  n_622;
assign n_625 = ~n_623 & ~n_624;
assign n_626 =  x_2276 & ~n_589;
assign n_627 =  i_26 &  n_589;
assign n_628 = ~n_626 & ~n_627;
assign n_629 =  x_2276 & ~n_628;
assign n_630 = ~x_2276 &  n_628;
assign n_631 = ~n_629 & ~n_630;
assign n_632 =  x_2275 & ~n_589;
assign n_633 =  i_25 &  n_589;
assign n_634 = ~n_632 & ~n_633;
assign n_635 =  x_2275 & ~n_634;
assign n_636 = ~x_2275 &  n_634;
assign n_637 = ~n_635 & ~n_636;
assign n_638 =  x_2274 & ~n_589;
assign n_639 =  i_24 &  n_589;
assign n_640 = ~n_638 & ~n_639;
assign n_641 =  x_2274 & ~n_640;
assign n_642 = ~x_2274 &  n_640;
assign n_643 = ~n_641 & ~n_642;
assign n_644 =  x_2273 & ~n_589;
assign n_645 =  i_23 &  n_589;
assign n_646 = ~n_644 & ~n_645;
assign n_647 =  x_2273 & ~n_646;
assign n_648 = ~x_2273 &  n_646;
assign n_649 = ~n_647 & ~n_648;
assign n_650 =  x_2272 & ~n_589;
assign n_651 =  i_22 &  n_589;
assign n_652 = ~n_650 & ~n_651;
assign n_653 =  x_2272 & ~n_652;
assign n_654 = ~x_2272 &  n_652;
assign n_655 = ~n_653 & ~n_654;
assign n_656 =  x_2271 & ~n_589;
assign n_657 =  i_21 &  n_589;
assign n_658 = ~n_656 & ~n_657;
assign n_659 =  x_2271 & ~n_658;
assign n_660 = ~x_2271 &  n_658;
assign n_661 = ~n_659 & ~n_660;
assign n_662 =  x_2270 & ~n_589;
assign n_663 =  i_20 &  n_589;
assign n_664 = ~n_662 & ~n_663;
assign n_665 =  x_2270 & ~n_664;
assign n_666 = ~x_2270 &  n_664;
assign n_667 = ~n_665 & ~n_666;
assign n_668 =  x_2269 & ~n_589;
assign n_669 =  i_19 &  n_589;
assign n_670 = ~n_668 & ~n_669;
assign n_671 =  x_2269 & ~n_670;
assign n_672 = ~x_2269 &  n_670;
assign n_673 = ~n_671 & ~n_672;
assign n_674 =  x_2268 & ~n_589;
assign n_675 =  i_18 &  n_589;
assign n_676 = ~n_674 & ~n_675;
assign n_677 =  x_2268 & ~n_676;
assign n_678 = ~x_2268 &  n_676;
assign n_679 = ~n_677 & ~n_678;
assign n_680 =  x_2267 & ~n_589;
assign n_681 =  i_17 &  n_589;
assign n_682 = ~n_680 & ~n_681;
assign n_683 =  x_2267 & ~n_682;
assign n_684 = ~x_2267 &  n_682;
assign n_685 = ~n_683 & ~n_684;
assign n_686 =  x_2266 & ~n_589;
assign n_687 =  i_16 &  n_589;
assign n_688 = ~n_686 & ~n_687;
assign n_689 =  x_2266 & ~n_688;
assign n_690 = ~x_2266 &  n_688;
assign n_691 = ~n_689 & ~n_690;
assign n_692 =  x_2265 & ~n_589;
assign n_693 =  i_15 &  n_589;
assign n_694 = ~n_692 & ~n_693;
assign n_695 =  x_2265 & ~n_694;
assign n_696 = ~x_2265 &  n_694;
assign n_697 = ~n_695 & ~n_696;
assign n_698 =  x_2264 & ~n_589;
assign n_699 =  i_14 &  n_589;
assign n_700 = ~n_698 & ~n_699;
assign n_701 =  x_2264 & ~n_700;
assign n_702 = ~x_2264 &  n_700;
assign n_703 = ~n_701 & ~n_702;
assign n_704 =  x_2263 & ~n_589;
assign n_705 =  i_13 &  n_589;
assign n_706 = ~n_704 & ~n_705;
assign n_707 =  x_2263 & ~n_706;
assign n_708 = ~x_2263 &  n_706;
assign n_709 = ~n_707 & ~n_708;
assign n_710 =  x_2262 & ~n_589;
assign n_711 =  i_12 &  n_589;
assign n_712 = ~n_710 & ~n_711;
assign n_713 =  x_2262 & ~n_712;
assign n_714 = ~x_2262 &  n_712;
assign n_715 = ~n_713 & ~n_714;
assign n_716 =  x_2261 & ~n_589;
assign n_717 =  i_11 &  n_589;
assign n_718 = ~n_716 & ~n_717;
assign n_719 =  x_2261 & ~n_718;
assign n_720 = ~x_2261 &  n_718;
assign n_721 = ~n_719 & ~n_720;
assign n_722 =  x_2260 & ~n_589;
assign n_723 =  i_10 &  n_589;
assign n_724 = ~n_722 & ~n_723;
assign n_725 =  x_2260 & ~n_724;
assign n_726 = ~x_2260 &  n_724;
assign n_727 = ~n_725 & ~n_726;
assign n_728 =  x_2259 & ~n_589;
assign n_729 =  i_9 &  n_589;
assign n_730 = ~n_728 & ~n_729;
assign n_731 =  x_2259 & ~n_730;
assign n_732 = ~x_2259 &  n_730;
assign n_733 = ~n_731 & ~n_732;
assign n_734 =  x_2258 & ~n_589;
assign n_735 =  i_8 &  n_589;
assign n_736 = ~n_734 & ~n_735;
assign n_737 =  x_2258 & ~n_736;
assign n_738 = ~x_2258 &  n_736;
assign n_739 = ~n_737 & ~n_738;
assign n_740 =  x_2257 & ~n_589;
assign n_741 =  i_7 &  n_589;
assign n_742 = ~n_740 & ~n_741;
assign n_743 =  x_2257 & ~n_742;
assign n_744 = ~x_2257 &  n_742;
assign n_745 = ~n_743 & ~n_744;
assign n_746 =  x_2256 & ~n_589;
assign n_747 =  i_6 &  n_589;
assign n_748 = ~n_746 & ~n_747;
assign n_749 =  x_2256 & ~n_748;
assign n_750 = ~x_2256 &  n_748;
assign n_751 = ~n_749 & ~n_750;
assign n_752 =  x_2255 & ~n_589;
assign n_753 =  i_5 &  n_589;
assign n_754 = ~n_752 & ~n_753;
assign n_755 =  x_2255 & ~n_754;
assign n_756 = ~x_2255 &  n_754;
assign n_757 = ~n_755 & ~n_756;
assign n_758 =  x_2254 & ~n_589;
assign n_759 =  i_4 &  n_589;
assign n_760 = ~n_758 & ~n_759;
assign n_761 =  x_2254 & ~n_760;
assign n_762 = ~x_2254 &  n_760;
assign n_763 = ~n_761 & ~n_762;
assign n_764 =  x_2253 & ~n_589;
assign n_765 =  i_3 &  n_589;
assign n_766 = ~n_764 & ~n_765;
assign n_767 =  x_2253 & ~n_766;
assign n_768 = ~x_2253 &  n_766;
assign n_769 = ~n_767 & ~n_768;
assign n_770 =  x_2252 & ~n_589;
assign n_771 =  i_2 &  n_589;
assign n_772 = ~n_770 & ~n_771;
assign n_773 =  x_2252 & ~n_772;
assign n_774 = ~x_2252 &  n_772;
assign n_775 = ~n_773 & ~n_774;
assign n_776 =  x_2251 & ~n_589;
assign n_777 =  i_1 &  n_589;
assign n_778 = ~n_776 & ~n_777;
assign n_779 =  x_2251 & ~n_778;
assign n_780 = ~x_2251 &  n_778;
assign n_781 = ~n_779 & ~n_780;
assign n_782 = ~x_39 &  x_40;
assign n_783 =  n_782 &  n_185;
assign n_784 = ~x_38 &  n_783;
assign n_785 = ~x_37 &  n_388;
assign n_786 =  n_784 &  n_785;
assign n_787 =  x_2250 & ~n_786;
assign n_788 =  i_32 &  n_786;
assign n_789 = ~n_787 & ~n_788;
assign n_790 =  x_2250 & ~n_789;
assign n_791 = ~x_2250 &  n_789;
assign n_792 = ~n_790 & ~n_791;
assign n_793 =  x_2249 & ~n_786;
assign n_794 =  i_31 &  n_786;
assign n_795 = ~n_793 & ~n_794;
assign n_796 =  x_2249 & ~n_795;
assign n_797 = ~x_2249 &  n_795;
assign n_798 = ~n_796 & ~n_797;
assign n_799 =  x_2248 & ~n_786;
assign n_800 =  i_30 &  n_786;
assign n_801 = ~n_799 & ~n_800;
assign n_802 =  x_2248 & ~n_801;
assign n_803 = ~x_2248 &  n_801;
assign n_804 = ~n_802 & ~n_803;
assign n_805 =  x_2247 & ~n_786;
assign n_806 =  i_29 &  n_786;
assign n_807 = ~n_805 & ~n_806;
assign n_808 =  x_2247 & ~n_807;
assign n_809 = ~x_2247 &  n_807;
assign n_810 = ~n_808 & ~n_809;
assign n_811 =  x_2246 & ~n_786;
assign n_812 =  i_28 &  n_786;
assign n_813 = ~n_811 & ~n_812;
assign n_814 =  x_2246 & ~n_813;
assign n_815 = ~x_2246 &  n_813;
assign n_816 = ~n_814 & ~n_815;
assign n_817 =  x_2245 & ~n_786;
assign n_818 =  i_27 &  n_786;
assign n_819 = ~n_817 & ~n_818;
assign n_820 =  x_2245 & ~n_819;
assign n_821 = ~x_2245 &  n_819;
assign n_822 = ~n_820 & ~n_821;
assign n_823 =  x_2244 & ~n_786;
assign n_824 =  i_26 &  n_786;
assign n_825 = ~n_823 & ~n_824;
assign n_826 =  x_2244 & ~n_825;
assign n_827 = ~x_2244 &  n_825;
assign n_828 = ~n_826 & ~n_827;
assign n_829 =  x_2243 & ~n_786;
assign n_830 =  i_25 &  n_786;
assign n_831 = ~n_829 & ~n_830;
assign n_832 =  x_2243 & ~n_831;
assign n_833 = ~x_2243 &  n_831;
assign n_834 = ~n_832 & ~n_833;
assign n_835 =  x_2242 & ~n_786;
assign n_836 =  i_24 &  n_786;
assign n_837 = ~n_835 & ~n_836;
assign n_838 =  x_2242 & ~n_837;
assign n_839 = ~x_2242 &  n_837;
assign n_840 = ~n_838 & ~n_839;
assign n_841 =  x_2241 & ~n_786;
assign n_842 =  i_23 &  n_786;
assign n_843 = ~n_841 & ~n_842;
assign n_844 =  x_2241 & ~n_843;
assign n_845 = ~x_2241 &  n_843;
assign n_846 = ~n_844 & ~n_845;
assign n_847 =  x_2240 & ~n_786;
assign n_848 =  i_22 &  n_786;
assign n_849 = ~n_847 & ~n_848;
assign n_850 =  x_2240 & ~n_849;
assign n_851 = ~x_2240 &  n_849;
assign n_852 = ~n_850 & ~n_851;
assign n_853 =  x_2239 & ~n_786;
assign n_854 =  i_21 &  n_786;
assign n_855 = ~n_853 & ~n_854;
assign n_856 =  x_2239 & ~n_855;
assign n_857 = ~x_2239 &  n_855;
assign n_858 = ~n_856 & ~n_857;
assign n_859 =  x_2238 & ~n_786;
assign n_860 =  i_20 &  n_786;
assign n_861 = ~n_859 & ~n_860;
assign n_862 =  x_2238 & ~n_861;
assign n_863 = ~x_2238 &  n_861;
assign n_864 = ~n_862 & ~n_863;
assign n_865 =  x_2237 & ~n_786;
assign n_866 =  i_19 &  n_786;
assign n_867 = ~n_865 & ~n_866;
assign n_868 =  x_2237 & ~n_867;
assign n_869 = ~x_2237 &  n_867;
assign n_870 = ~n_868 & ~n_869;
assign n_871 =  x_2236 & ~n_786;
assign n_872 =  i_18 &  n_786;
assign n_873 = ~n_871 & ~n_872;
assign n_874 =  x_2236 & ~n_873;
assign n_875 = ~x_2236 &  n_873;
assign n_876 = ~n_874 & ~n_875;
assign n_877 =  x_2235 & ~n_786;
assign n_878 =  i_17 &  n_786;
assign n_879 = ~n_877 & ~n_878;
assign n_880 =  x_2235 & ~n_879;
assign n_881 = ~x_2235 &  n_879;
assign n_882 = ~n_880 & ~n_881;
assign n_883 =  x_2234 & ~n_786;
assign n_884 =  i_16 &  n_786;
assign n_885 = ~n_883 & ~n_884;
assign n_886 =  x_2234 & ~n_885;
assign n_887 = ~x_2234 &  n_885;
assign n_888 = ~n_886 & ~n_887;
assign n_889 =  x_2233 & ~n_786;
assign n_890 =  i_15 &  n_786;
assign n_891 = ~n_889 & ~n_890;
assign n_892 =  x_2233 & ~n_891;
assign n_893 = ~x_2233 &  n_891;
assign n_894 = ~n_892 & ~n_893;
assign n_895 =  x_2232 & ~n_786;
assign n_896 =  i_14 &  n_786;
assign n_897 = ~n_895 & ~n_896;
assign n_898 =  x_2232 & ~n_897;
assign n_899 = ~x_2232 &  n_897;
assign n_900 = ~n_898 & ~n_899;
assign n_901 =  x_2231 & ~n_786;
assign n_902 =  i_13 &  n_786;
assign n_903 = ~n_901 & ~n_902;
assign n_904 =  x_2231 & ~n_903;
assign n_905 = ~x_2231 &  n_903;
assign n_906 = ~n_904 & ~n_905;
assign n_907 =  x_2230 & ~n_786;
assign n_908 =  i_12 &  n_786;
assign n_909 = ~n_907 & ~n_908;
assign n_910 =  x_2230 & ~n_909;
assign n_911 = ~x_2230 &  n_909;
assign n_912 = ~n_910 & ~n_911;
assign n_913 =  x_2229 & ~n_786;
assign n_914 =  i_11 &  n_786;
assign n_915 = ~n_913 & ~n_914;
assign n_916 =  x_2229 & ~n_915;
assign n_917 = ~x_2229 &  n_915;
assign n_918 = ~n_916 & ~n_917;
assign n_919 =  x_2228 & ~n_786;
assign n_920 =  i_10 &  n_786;
assign n_921 = ~n_919 & ~n_920;
assign n_922 =  x_2228 & ~n_921;
assign n_923 = ~x_2228 &  n_921;
assign n_924 = ~n_922 & ~n_923;
assign n_925 =  x_2227 & ~n_786;
assign n_926 =  i_9 &  n_786;
assign n_927 = ~n_925 & ~n_926;
assign n_928 =  x_2227 & ~n_927;
assign n_929 = ~x_2227 &  n_927;
assign n_930 = ~n_928 & ~n_929;
assign n_931 =  x_2226 & ~n_786;
assign n_932 =  i_8 &  n_786;
assign n_933 = ~n_931 & ~n_932;
assign n_934 =  x_2226 & ~n_933;
assign n_935 = ~x_2226 &  n_933;
assign n_936 = ~n_934 & ~n_935;
assign n_937 =  x_2225 & ~n_786;
assign n_938 =  i_7 &  n_786;
assign n_939 = ~n_937 & ~n_938;
assign n_940 =  x_2225 & ~n_939;
assign n_941 = ~x_2225 &  n_939;
assign n_942 = ~n_940 & ~n_941;
assign n_943 =  x_2224 & ~n_786;
assign n_944 =  i_6 &  n_786;
assign n_945 = ~n_943 & ~n_944;
assign n_946 =  x_2224 & ~n_945;
assign n_947 = ~x_2224 &  n_945;
assign n_948 = ~n_946 & ~n_947;
assign n_949 =  x_2223 & ~n_786;
assign n_950 =  i_5 &  n_786;
assign n_951 = ~n_949 & ~n_950;
assign n_952 =  x_2223 & ~n_951;
assign n_953 = ~x_2223 &  n_951;
assign n_954 = ~n_952 & ~n_953;
assign n_955 =  x_2222 & ~n_786;
assign n_956 =  i_4 &  n_786;
assign n_957 = ~n_955 & ~n_956;
assign n_958 =  x_2222 & ~n_957;
assign n_959 = ~x_2222 &  n_957;
assign n_960 = ~n_958 & ~n_959;
assign n_961 =  x_2221 & ~n_786;
assign n_962 =  i_3 &  n_786;
assign n_963 = ~n_961 & ~n_962;
assign n_964 =  x_2221 & ~n_963;
assign n_965 = ~x_2221 &  n_963;
assign n_966 = ~n_964 & ~n_965;
assign n_967 =  x_2220 & ~n_786;
assign n_968 =  i_2 &  n_786;
assign n_969 = ~n_967 & ~n_968;
assign n_970 =  x_2220 & ~n_969;
assign n_971 = ~x_2220 &  n_969;
assign n_972 = ~n_970 & ~n_971;
assign n_973 =  x_2219 & ~n_786;
assign n_974 =  i_1 &  n_786;
assign n_975 = ~n_973 & ~n_974;
assign n_976 =  x_2219 & ~n_975;
assign n_977 = ~x_2219 &  n_975;
assign n_978 = ~n_976 & ~n_977;
assign n_979 = ~x_41 &  x_42;
assign n_980 =  n_184 &  n_979;
assign n_981 =  x_35 &  n_189;
assign n_982 =  x_36 &  n_981;
assign n_983 =  n_4 &  n_982;
assign n_984 =  n_980 &  n_983;
assign n_985 =  i_32 &  n_984;
assign n_986 =  x_2218 & ~n_984;
assign n_987 = ~n_985 & ~n_986;
assign n_988 =  x_2218 & ~n_987;
assign n_989 = ~x_2218 &  n_987;
assign n_990 = ~n_988 & ~n_989;
assign n_991 =  i_31 &  n_984;
assign n_992 =  x_2217 & ~n_984;
assign n_993 = ~n_991 & ~n_992;
assign n_994 =  x_2217 & ~n_993;
assign n_995 = ~x_2217 &  n_993;
assign n_996 = ~n_994 & ~n_995;
assign n_997 =  i_30 &  n_984;
assign n_998 =  x_2216 & ~n_984;
assign n_999 = ~n_997 & ~n_998;
assign n_1000 =  x_2216 & ~n_999;
assign n_1001 = ~x_2216 &  n_999;
assign n_1002 = ~n_1000 & ~n_1001;
assign n_1003 =  i_29 &  n_984;
assign n_1004 =  x_2215 & ~n_984;
assign n_1005 = ~n_1003 & ~n_1004;
assign n_1006 =  x_2215 & ~n_1005;
assign n_1007 = ~x_2215 &  n_1005;
assign n_1008 = ~n_1006 & ~n_1007;
assign n_1009 =  i_28 &  n_984;
assign n_1010 =  x_2214 & ~n_984;
assign n_1011 = ~n_1009 & ~n_1010;
assign n_1012 =  x_2214 & ~n_1011;
assign n_1013 = ~x_2214 &  n_1011;
assign n_1014 = ~n_1012 & ~n_1013;
assign n_1015 =  i_27 &  n_984;
assign n_1016 =  x_2213 & ~n_984;
assign n_1017 = ~n_1015 & ~n_1016;
assign n_1018 =  x_2213 & ~n_1017;
assign n_1019 = ~x_2213 &  n_1017;
assign n_1020 = ~n_1018 & ~n_1019;
assign n_1021 =  i_26 &  n_984;
assign n_1022 =  x_2212 & ~n_984;
assign n_1023 = ~n_1021 & ~n_1022;
assign n_1024 =  x_2212 & ~n_1023;
assign n_1025 = ~x_2212 &  n_1023;
assign n_1026 = ~n_1024 & ~n_1025;
assign n_1027 =  i_25 &  n_984;
assign n_1028 =  x_2211 & ~n_984;
assign n_1029 = ~n_1027 & ~n_1028;
assign n_1030 =  x_2211 & ~n_1029;
assign n_1031 = ~x_2211 &  n_1029;
assign n_1032 = ~n_1030 & ~n_1031;
assign n_1033 =  i_24 &  n_984;
assign n_1034 =  x_2210 & ~n_984;
assign n_1035 = ~n_1033 & ~n_1034;
assign n_1036 =  x_2210 & ~n_1035;
assign n_1037 = ~x_2210 &  n_1035;
assign n_1038 = ~n_1036 & ~n_1037;
assign n_1039 =  i_23 &  n_984;
assign n_1040 =  x_2209 & ~n_984;
assign n_1041 = ~n_1039 & ~n_1040;
assign n_1042 =  x_2209 & ~n_1041;
assign n_1043 = ~x_2209 &  n_1041;
assign n_1044 = ~n_1042 & ~n_1043;
assign n_1045 =  i_22 &  n_984;
assign n_1046 =  x_2208 & ~n_984;
assign n_1047 = ~n_1045 & ~n_1046;
assign n_1048 =  x_2208 & ~n_1047;
assign n_1049 = ~x_2208 &  n_1047;
assign n_1050 = ~n_1048 & ~n_1049;
assign n_1051 =  i_21 &  n_984;
assign n_1052 =  x_2207 & ~n_984;
assign n_1053 = ~n_1051 & ~n_1052;
assign n_1054 =  x_2207 & ~n_1053;
assign n_1055 = ~x_2207 &  n_1053;
assign n_1056 = ~n_1054 & ~n_1055;
assign n_1057 =  i_20 &  n_984;
assign n_1058 =  x_2206 & ~n_984;
assign n_1059 = ~n_1057 & ~n_1058;
assign n_1060 =  x_2206 & ~n_1059;
assign n_1061 = ~x_2206 &  n_1059;
assign n_1062 = ~n_1060 & ~n_1061;
assign n_1063 =  i_19 &  n_984;
assign n_1064 =  x_2205 & ~n_984;
assign n_1065 = ~n_1063 & ~n_1064;
assign n_1066 =  x_2205 & ~n_1065;
assign n_1067 = ~x_2205 &  n_1065;
assign n_1068 = ~n_1066 & ~n_1067;
assign n_1069 =  i_18 &  n_984;
assign n_1070 =  x_2204 & ~n_984;
assign n_1071 = ~n_1069 & ~n_1070;
assign n_1072 =  x_2204 & ~n_1071;
assign n_1073 = ~x_2204 &  n_1071;
assign n_1074 = ~n_1072 & ~n_1073;
assign n_1075 =  i_17 &  n_984;
assign n_1076 =  x_2203 & ~n_984;
assign n_1077 = ~n_1075 & ~n_1076;
assign n_1078 =  x_2203 & ~n_1077;
assign n_1079 = ~x_2203 &  n_1077;
assign n_1080 = ~n_1078 & ~n_1079;
assign n_1081 =  i_16 &  n_984;
assign n_1082 =  x_2202 & ~n_984;
assign n_1083 = ~n_1081 & ~n_1082;
assign n_1084 =  x_2202 & ~n_1083;
assign n_1085 = ~x_2202 &  n_1083;
assign n_1086 = ~n_1084 & ~n_1085;
assign n_1087 =  i_15 &  n_984;
assign n_1088 =  x_2201 & ~n_984;
assign n_1089 = ~n_1087 & ~n_1088;
assign n_1090 =  x_2201 & ~n_1089;
assign n_1091 = ~x_2201 &  n_1089;
assign n_1092 = ~n_1090 & ~n_1091;
assign n_1093 =  i_14 &  n_984;
assign n_1094 =  x_2200 & ~n_984;
assign n_1095 = ~n_1093 & ~n_1094;
assign n_1096 =  x_2200 & ~n_1095;
assign n_1097 = ~x_2200 &  n_1095;
assign n_1098 = ~n_1096 & ~n_1097;
assign n_1099 =  i_13 &  n_984;
assign n_1100 =  x_2199 & ~n_984;
assign n_1101 = ~n_1099 & ~n_1100;
assign n_1102 =  x_2199 & ~n_1101;
assign n_1103 = ~x_2199 &  n_1101;
assign n_1104 = ~n_1102 & ~n_1103;
assign n_1105 =  i_12 &  n_984;
assign n_1106 =  x_2198 & ~n_984;
assign n_1107 = ~n_1105 & ~n_1106;
assign n_1108 =  x_2198 & ~n_1107;
assign n_1109 = ~x_2198 &  n_1107;
assign n_1110 = ~n_1108 & ~n_1109;
assign n_1111 =  i_11 &  n_984;
assign n_1112 =  x_2197 & ~n_984;
assign n_1113 = ~n_1111 & ~n_1112;
assign n_1114 =  x_2197 & ~n_1113;
assign n_1115 = ~x_2197 &  n_1113;
assign n_1116 = ~n_1114 & ~n_1115;
assign n_1117 =  i_10 &  n_984;
assign n_1118 =  x_2196 & ~n_984;
assign n_1119 = ~n_1117 & ~n_1118;
assign n_1120 =  x_2196 & ~n_1119;
assign n_1121 = ~x_2196 &  n_1119;
assign n_1122 = ~n_1120 & ~n_1121;
assign n_1123 =  i_9 &  n_984;
assign n_1124 =  x_2195 & ~n_984;
assign n_1125 = ~n_1123 & ~n_1124;
assign n_1126 =  x_2195 & ~n_1125;
assign n_1127 = ~x_2195 &  n_1125;
assign n_1128 = ~n_1126 & ~n_1127;
assign n_1129 =  i_8 &  n_984;
assign n_1130 =  x_2194 & ~n_984;
assign n_1131 = ~n_1129 & ~n_1130;
assign n_1132 =  x_2194 & ~n_1131;
assign n_1133 = ~x_2194 &  n_1131;
assign n_1134 = ~n_1132 & ~n_1133;
assign n_1135 =  i_7 &  n_984;
assign n_1136 =  x_2193 & ~n_984;
assign n_1137 = ~n_1135 & ~n_1136;
assign n_1138 =  x_2193 & ~n_1137;
assign n_1139 = ~x_2193 &  n_1137;
assign n_1140 = ~n_1138 & ~n_1139;
assign n_1141 =  i_6 &  n_984;
assign n_1142 =  x_2192 & ~n_984;
assign n_1143 = ~n_1141 & ~n_1142;
assign n_1144 =  x_2192 & ~n_1143;
assign n_1145 = ~x_2192 &  n_1143;
assign n_1146 = ~n_1144 & ~n_1145;
assign n_1147 =  i_5 &  n_984;
assign n_1148 =  x_2191 & ~n_984;
assign n_1149 = ~n_1147 & ~n_1148;
assign n_1150 =  x_2191 & ~n_1149;
assign n_1151 = ~x_2191 &  n_1149;
assign n_1152 = ~n_1150 & ~n_1151;
assign n_1153 =  i_4 &  n_984;
assign n_1154 =  x_2190 & ~n_984;
assign n_1155 = ~n_1153 & ~n_1154;
assign n_1156 =  x_2190 & ~n_1155;
assign n_1157 = ~x_2190 &  n_1155;
assign n_1158 = ~n_1156 & ~n_1157;
assign n_1159 =  i_3 &  n_984;
assign n_1160 =  x_2189 & ~n_984;
assign n_1161 = ~n_1159 & ~n_1160;
assign n_1162 =  x_2189 & ~n_1161;
assign n_1163 = ~x_2189 &  n_1161;
assign n_1164 = ~n_1162 & ~n_1163;
assign n_1165 =  i_2 &  n_984;
assign n_1166 =  x_2188 & ~n_984;
assign n_1167 = ~n_1165 & ~n_1166;
assign n_1168 =  x_2188 & ~n_1167;
assign n_1169 = ~x_2188 &  n_1167;
assign n_1170 = ~n_1168 & ~n_1169;
assign n_1171 =  i_1 &  n_984;
assign n_1172 =  x_2187 & ~n_984;
assign n_1173 = ~n_1171 & ~n_1172;
assign n_1174 =  x_2187 & ~n_1173;
assign n_1175 = ~x_2187 &  n_1173;
assign n_1176 = ~n_1174 & ~n_1175;
assign n_1177 = ~x_35 & ~x_36;
assign n_1178 =  n_189 &  n_1177;
assign n_1179 =  n_4 &  n_1178;
assign n_1180 =  n_385 &  n_1179;
assign n_1181 =  x_42 &  n_1180;
assign n_1182 =  x_2186 & ~n_1180;
assign n_1183 = ~n_1181 & ~n_1182;
assign n_1184 =  x_2186 & ~n_1183;
assign n_1185 = ~x_2186 &  n_1183;
assign n_1186 = ~n_1184 & ~n_1185;
assign n_1187 =  x_2185 & ~n_1180;
assign n_1188 =  x_2185 &  n_1187;
assign n_1189 = ~x_2185 & ~n_1187;
assign n_1190 = ~n_1188 & ~n_1189;
assign n_1191 =  x_2184 & ~n_1180;
assign n_1192 =  x_2184 &  n_1191;
assign n_1193 = ~x_2184 & ~n_1191;
assign n_1194 = ~n_1192 & ~n_1193;
assign n_1195 =  x_2183 & ~n_1180;
assign n_1196 =  x_2183 &  n_1195;
assign n_1197 = ~x_2183 & ~n_1195;
assign n_1198 = ~n_1196 & ~n_1197;
assign n_1199 =  x_2182 & ~n_1180;
assign n_1200 =  x_2182 &  n_1199;
assign n_1201 = ~x_2182 & ~n_1199;
assign n_1202 = ~n_1200 & ~n_1201;
assign n_1203 =  x_2181 & ~n_1180;
assign n_1204 =  x_2181 &  n_1203;
assign n_1205 = ~x_2181 & ~n_1203;
assign n_1206 = ~n_1204 & ~n_1205;
assign n_1207 =  x_2180 & ~n_1180;
assign n_1208 =  x_2180 &  n_1207;
assign n_1209 = ~x_2180 & ~n_1207;
assign n_1210 = ~n_1208 & ~n_1209;
assign n_1211 =  x_2179 & ~n_1180;
assign n_1212 =  x_2179 &  n_1211;
assign n_1213 = ~x_2179 & ~n_1211;
assign n_1214 = ~n_1212 & ~n_1213;
assign n_1215 =  x_2178 & ~n_1180;
assign n_1216 =  x_2178 &  n_1215;
assign n_1217 = ~x_2178 & ~n_1215;
assign n_1218 = ~n_1216 & ~n_1217;
assign n_1219 =  x_2177 & ~n_1180;
assign n_1220 =  x_2177 &  n_1219;
assign n_1221 = ~x_2177 & ~n_1219;
assign n_1222 = ~n_1220 & ~n_1221;
assign n_1223 =  x_2176 & ~n_1180;
assign n_1224 =  x_2176 &  n_1223;
assign n_1225 = ~x_2176 & ~n_1223;
assign n_1226 = ~n_1224 & ~n_1225;
assign n_1227 =  x_2175 & ~n_1180;
assign n_1228 =  x_2175 &  n_1227;
assign n_1229 = ~x_2175 & ~n_1227;
assign n_1230 = ~n_1228 & ~n_1229;
assign n_1231 =  x_2174 & ~n_1180;
assign n_1232 =  x_2174 &  n_1231;
assign n_1233 = ~x_2174 & ~n_1231;
assign n_1234 = ~n_1232 & ~n_1233;
assign n_1235 =  x_2173 & ~n_1180;
assign n_1236 =  x_2173 &  n_1235;
assign n_1237 = ~x_2173 & ~n_1235;
assign n_1238 = ~n_1236 & ~n_1237;
assign n_1239 =  x_2172 & ~n_1180;
assign n_1240 =  x_2172 &  n_1239;
assign n_1241 = ~x_2172 & ~n_1239;
assign n_1242 = ~n_1240 & ~n_1241;
assign n_1243 =  x_2171 & ~n_1180;
assign n_1244 =  x_2171 &  n_1243;
assign n_1245 = ~x_2171 & ~n_1243;
assign n_1246 = ~n_1244 & ~n_1245;
assign n_1247 =  x_2170 & ~n_1180;
assign n_1248 =  x_2170 &  n_1247;
assign n_1249 = ~x_2170 & ~n_1247;
assign n_1250 = ~n_1248 & ~n_1249;
assign n_1251 =  x_2169 & ~n_1180;
assign n_1252 =  x_2169 &  n_1251;
assign n_1253 = ~x_2169 & ~n_1251;
assign n_1254 = ~n_1252 & ~n_1253;
assign n_1255 =  x_2168 & ~n_1180;
assign n_1256 =  x_2168 &  n_1255;
assign n_1257 = ~x_2168 & ~n_1255;
assign n_1258 = ~n_1256 & ~n_1257;
assign n_1259 =  x_2167 & ~n_1180;
assign n_1260 =  x_2167 &  n_1259;
assign n_1261 = ~x_2167 & ~n_1259;
assign n_1262 = ~n_1260 & ~n_1261;
assign n_1263 =  x_2166 & ~n_1180;
assign n_1264 =  x_2166 &  n_1263;
assign n_1265 = ~x_2166 & ~n_1263;
assign n_1266 = ~n_1264 & ~n_1265;
assign n_1267 =  x_2165 & ~n_1180;
assign n_1268 =  x_2165 &  n_1267;
assign n_1269 = ~x_2165 & ~n_1267;
assign n_1270 = ~n_1268 & ~n_1269;
assign n_1271 =  x_2164 & ~n_1180;
assign n_1272 =  x_2164 &  n_1271;
assign n_1273 = ~x_2164 & ~n_1271;
assign n_1274 = ~n_1272 & ~n_1273;
assign n_1275 =  x_2163 & ~n_1180;
assign n_1276 =  x_2163 &  n_1275;
assign n_1277 = ~x_2163 & ~n_1275;
assign n_1278 = ~n_1276 & ~n_1277;
assign n_1279 =  x_2162 & ~n_1180;
assign n_1280 =  x_2162 &  n_1279;
assign n_1281 = ~x_2162 & ~n_1279;
assign n_1282 = ~n_1280 & ~n_1281;
assign n_1283 =  x_2161 & ~n_1180;
assign n_1284 =  x_2161 &  n_1283;
assign n_1285 = ~x_2161 & ~n_1283;
assign n_1286 = ~n_1284 & ~n_1285;
assign n_1287 =  x_2160 & ~n_1180;
assign n_1288 =  x_2160 &  n_1287;
assign n_1289 = ~x_2160 & ~n_1287;
assign n_1290 = ~n_1288 & ~n_1289;
assign n_1291 =  x_2159 & ~n_1180;
assign n_1292 =  x_2159 &  n_1291;
assign n_1293 = ~x_2159 & ~n_1291;
assign n_1294 = ~n_1292 & ~n_1293;
assign n_1295 =  x_2158 & ~n_1180;
assign n_1296 =  x_2158 &  n_1295;
assign n_1297 = ~x_2158 & ~n_1295;
assign n_1298 = ~n_1296 & ~n_1297;
assign n_1299 =  x_2157 & ~n_1180;
assign n_1300 =  x_2157 &  n_1299;
assign n_1301 = ~x_2157 & ~n_1299;
assign n_1302 = ~n_1300 & ~n_1301;
assign n_1303 =  x_2156 & ~n_1180;
assign n_1304 =  x_2156 &  n_1303;
assign n_1305 = ~x_2156 & ~n_1303;
assign n_1306 = ~n_1304 & ~n_1305;
assign n_1307 =  x_2155 & ~n_1180;
assign n_1308 =  x_2155 &  n_1307;
assign n_1309 = ~x_2155 & ~n_1307;
assign n_1310 = ~n_1308 & ~n_1309;
assign n_1311 =  x_36 & ~x_37;
assign n_1312 = ~x_38 &  n_1311;
assign n_1313 = ~x_39 &  n_1312;
assign n_1314 = ~x_40 & ~x_41;
assign n_1315 = ~x_42 &  n_1314;
assign n_1316 =  n_387 &  n_1315;
assign n_1317 =  n_1313 &  n_1316;
assign n_1318 =  x_2154 & ~n_1317;
assign n_1319 =  i_32 &  n_1317;
assign n_1320 = ~n_1318 & ~n_1319;
assign n_1321 =  x_2154 & ~n_1320;
assign n_1322 = ~x_2154 &  n_1320;
assign n_1323 = ~n_1321 & ~n_1322;
assign n_1324 =  x_2153 & ~n_1317;
assign n_1325 =  i_31 &  n_1317;
assign n_1326 = ~n_1324 & ~n_1325;
assign n_1327 =  x_2153 & ~n_1326;
assign n_1328 = ~x_2153 &  n_1326;
assign n_1329 = ~n_1327 & ~n_1328;
assign n_1330 =  x_2152 & ~n_1317;
assign n_1331 =  i_30 &  n_1317;
assign n_1332 = ~n_1330 & ~n_1331;
assign n_1333 =  x_2152 & ~n_1332;
assign n_1334 = ~x_2152 &  n_1332;
assign n_1335 = ~n_1333 & ~n_1334;
assign n_1336 =  x_2151 & ~n_1317;
assign n_1337 =  i_29 &  n_1317;
assign n_1338 = ~n_1336 & ~n_1337;
assign n_1339 =  x_2151 & ~n_1338;
assign n_1340 = ~x_2151 &  n_1338;
assign n_1341 = ~n_1339 & ~n_1340;
assign n_1342 =  x_2150 & ~n_1317;
assign n_1343 =  i_28 &  n_1317;
assign n_1344 = ~n_1342 & ~n_1343;
assign n_1345 =  x_2150 & ~n_1344;
assign n_1346 = ~x_2150 &  n_1344;
assign n_1347 = ~n_1345 & ~n_1346;
assign n_1348 =  x_2149 & ~n_1317;
assign n_1349 =  i_27 &  n_1317;
assign n_1350 = ~n_1348 & ~n_1349;
assign n_1351 =  x_2149 & ~n_1350;
assign n_1352 = ~x_2149 &  n_1350;
assign n_1353 = ~n_1351 & ~n_1352;
assign n_1354 =  x_2148 & ~n_1317;
assign n_1355 =  i_26 &  n_1317;
assign n_1356 = ~n_1354 & ~n_1355;
assign n_1357 =  x_2148 & ~n_1356;
assign n_1358 = ~x_2148 &  n_1356;
assign n_1359 = ~n_1357 & ~n_1358;
assign n_1360 =  x_2147 & ~n_1317;
assign n_1361 =  i_25 &  n_1317;
assign n_1362 = ~n_1360 & ~n_1361;
assign n_1363 =  x_2147 & ~n_1362;
assign n_1364 = ~x_2147 &  n_1362;
assign n_1365 = ~n_1363 & ~n_1364;
assign n_1366 =  x_2146 & ~n_1317;
assign n_1367 =  i_24 &  n_1317;
assign n_1368 = ~n_1366 & ~n_1367;
assign n_1369 =  x_2146 & ~n_1368;
assign n_1370 = ~x_2146 &  n_1368;
assign n_1371 = ~n_1369 & ~n_1370;
assign n_1372 =  x_2145 & ~n_1317;
assign n_1373 =  i_23 &  n_1317;
assign n_1374 = ~n_1372 & ~n_1373;
assign n_1375 =  x_2145 & ~n_1374;
assign n_1376 = ~x_2145 &  n_1374;
assign n_1377 = ~n_1375 & ~n_1376;
assign n_1378 =  x_2144 & ~n_1317;
assign n_1379 =  i_22 &  n_1317;
assign n_1380 = ~n_1378 & ~n_1379;
assign n_1381 =  x_2144 & ~n_1380;
assign n_1382 = ~x_2144 &  n_1380;
assign n_1383 = ~n_1381 & ~n_1382;
assign n_1384 =  x_2143 & ~n_1317;
assign n_1385 =  i_21 &  n_1317;
assign n_1386 = ~n_1384 & ~n_1385;
assign n_1387 =  x_2143 & ~n_1386;
assign n_1388 = ~x_2143 &  n_1386;
assign n_1389 = ~n_1387 & ~n_1388;
assign n_1390 =  x_2142 & ~n_1317;
assign n_1391 =  i_20 &  n_1317;
assign n_1392 = ~n_1390 & ~n_1391;
assign n_1393 =  x_2142 & ~n_1392;
assign n_1394 = ~x_2142 &  n_1392;
assign n_1395 = ~n_1393 & ~n_1394;
assign n_1396 =  x_2141 & ~n_1317;
assign n_1397 =  i_19 &  n_1317;
assign n_1398 = ~n_1396 & ~n_1397;
assign n_1399 =  x_2141 & ~n_1398;
assign n_1400 = ~x_2141 &  n_1398;
assign n_1401 = ~n_1399 & ~n_1400;
assign n_1402 =  x_2140 & ~n_1317;
assign n_1403 =  i_18 &  n_1317;
assign n_1404 = ~n_1402 & ~n_1403;
assign n_1405 =  x_2140 & ~n_1404;
assign n_1406 = ~x_2140 &  n_1404;
assign n_1407 = ~n_1405 & ~n_1406;
assign n_1408 =  x_2139 & ~n_1317;
assign n_1409 =  i_17 &  n_1317;
assign n_1410 = ~n_1408 & ~n_1409;
assign n_1411 =  x_2139 & ~n_1410;
assign n_1412 = ~x_2139 &  n_1410;
assign n_1413 = ~n_1411 & ~n_1412;
assign n_1414 =  x_2138 & ~n_1317;
assign n_1415 =  i_16 &  n_1317;
assign n_1416 = ~n_1414 & ~n_1415;
assign n_1417 =  x_2138 & ~n_1416;
assign n_1418 = ~x_2138 &  n_1416;
assign n_1419 = ~n_1417 & ~n_1418;
assign n_1420 =  x_2137 & ~n_1317;
assign n_1421 =  i_15 &  n_1317;
assign n_1422 = ~n_1420 & ~n_1421;
assign n_1423 =  x_2137 & ~n_1422;
assign n_1424 = ~x_2137 &  n_1422;
assign n_1425 = ~n_1423 & ~n_1424;
assign n_1426 =  x_2136 & ~n_1317;
assign n_1427 =  i_14 &  n_1317;
assign n_1428 = ~n_1426 & ~n_1427;
assign n_1429 =  x_2136 & ~n_1428;
assign n_1430 = ~x_2136 &  n_1428;
assign n_1431 = ~n_1429 & ~n_1430;
assign n_1432 =  x_2135 & ~n_1317;
assign n_1433 =  i_13 &  n_1317;
assign n_1434 = ~n_1432 & ~n_1433;
assign n_1435 =  x_2135 & ~n_1434;
assign n_1436 = ~x_2135 &  n_1434;
assign n_1437 = ~n_1435 & ~n_1436;
assign n_1438 =  x_2134 & ~n_1317;
assign n_1439 =  i_12 &  n_1317;
assign n_1440 = ~n_1438 & ~n_1439;
assign n_1441 =  x_2134 & ~n_1440;
assign n_1442 = ~x_2134 &  n_1440;
assign n_1443 = ~n_1441 & ~n_1442;
assign n_1444 =  x_2133 & ~n_1317;
assign n_1445 =  i_11 &  n_1317;
assign n_1446 = ~n_1444 & ~n_1445;
assign n_1447 =  x_2133 & ~n_1446;
assign n_1448 = ~x_2133 &  n_1446;
assign n_1449 = ~n_1447 & ~n_1448;
assign n_1450 =  x_2132 & ~n_1317;
assign n_1451 =  i_10 &  n_1317;
assign n_1452 = ~n_1450 & ~n_1451;
assign n_1453 =  x_2132 & ~n_1452;
assign n_1454 = ~x_2132 &  n_1452;
assign n_1455 = ~n_1453 & ~n_1454;
assign n_1456 =  x_2131 & ~n_1317;
assign n_1457 =  i_9 &  n_1317;
assign n_1458 = ~n_1456 & ~n_1457;
assign n_1459 =  x_2131 & ~n_1458;
assign n_1460 = ~x_2131 &  n_1458;
assign n_1461 = ~n_1459 & ~n_1460;
assign n_1462 =  x_2130 & ~n_1317;
assign n_1463 =  i_8 &  n_1317;
assign n_1464 = ~n_1462 & ~n_1463;
assign n_1465 =  x_2130 & ~n_1464;
assign n_1466 = ~x_2130 &  n_1464;
assign n_1467 = ~n_1465 & ~n_1466;
assign n_1468 =  x_2129 & ~n_1317;
assign n_1469 =  i_7 &  n_1317;
assign n_1470 = ~n_1468 & ~n_1469;
assign n_1471 =  x_2129 & ~n_1470;
assign n_1472 = ~x_2129 &  n_1470;
assign n_1473 = ~n_1471 & ~n_1472;
assign n_1474 =  x_2128 & ~n_1317;
assign n_1475 =  i_6 &  n_1317;
assign n_1476 = ~n_1474 & ~n_1475;
assign n_1477 =  x_2128 & ~n_1476;
assign n_1478 = ~x_2128 &  n_1476;
assign n_1479 = ~n_1477 & ~n_1478;
assign n_1480 =  x_2127 & ~n_1317;
assign n_1481 =  i_5 &  n_1317;
assign n_1482 = ~n_1480 & ~n_1481;
assign n_1483 =  x_2127 & ~n_1482;
assign n_1484 = ~x_2127 &  n_1482;
assign n_1485 = ~n_1483 & ~n_1484;
assign n_1486 =  x_2126 & ~n_1317;
assign n_1487 =  i_4 &  n_1317;
assign n_1488 = ~n_1486 & ~n_1487;
assign n_1489 =  x_2126 & ~n_1488;
assign n_1490 = ~x_2126 &  n_1488;
assign n_1491 = ~n_1489 & ~n_1490;
assign n_1492 =  x_2125 & ~n_1317;
assign n_1493 =  i_3 &  n_1317;
assign n_1494 = ~n_1492 & ~n_1493;
assign n_1495 =  x_2125 & ~n_1494;
assign n_1496 = ~x_2125 &  n_1494;
assign n_1497 = ~n_1495 & ~n_1496;
assign n_1498 =  x_2124 & ~n_1317;
assign n_1499 =  i_2 &  n_1317;
assign n_1500 = ~n_1498 & ~n_1499;
assign n_1501 =  x_2124 & ~n_1500;
assign n_1502 = ~x_2124 &  n_1500;
assign n_1503 = ~n_1501 & ~n_1502;
assign n_1504 =  x_2123 & ~n_1317;
assign n_1505 =  i_1 &  n_1317;
assign n_1506 = ~n_1504 & ~n_1505;
assign n_1507 =  x_2123 & ~n_1506;
assign n_1508 = ~x_2123 &  n_1506;
assign n_1509 = ~n_1507 & ~n_1508;
assign n_1510 = ~x_38 &  x_39;
assign n_1511 = ~x_37 &  n_190;
assign n_1512 =  n_1510 &  n_1511;
assign n_1513 =  n_1512 &  n_2;
assign n_1514 =  x_2122 & ~n_1513;
assign n_1515 =  i_32 &  n_1513;
assign n_1516 = ~n_1514 & ~n_1515;
assign n_1517 =  x_2122 & ~n_1516;
assign n_1518 = ~x_2122 &  n_1516;
assign n_1519 = ~n_1517 & ~n_1518;
assign n_1520 =  x_2121 & ~n_1513;
assign n_1521 =  i_31 &  n_1513;
assign n_1522 = ~n_1520 & ~n_1521;
assign n_1523 =  x_2121 & ~n_1522;
assign n_1524 = ~x_2121 &  n_1522;
assign n_1525 = ~n_1523 & ~n_1524;
assign n_1526 =  x_2120 & ~n_1513;
assign n_1527 =  i_30 &  n_1513;
assign n_1528 = ~n_1526 & ~n_1527;
assign n_1529 =  x_2120 & ~n_1528;
assign n_1530 = ~x_2120 &  n_1528;
assign n_1531 = ~n_1529 & ~n_1530;
assign n_1532 =  x_2119 & ~n_1513;
assign n_1533 =  i_29 &  n_1513;
assign n_1534 = ~n_1532 & ~n_1533;
assign n_1535 =  x_2119 & ~n_1534;
assign n_1536 = ~x_2119 &  n_1534;
assign n_1537 = ~n_1535 & ~n_1536;
assign n_1538 =  x_2118 & ~n_1513;
assign n_1539 =  i_28 &  n_1513;
assign n_1540 = ~n_1538 & ~n_1539;
assign n_1541 =  x_2118 & ~n_1540;
assign n_1542 = ~x_2118 &  n_1540;
assign n_1543 = ~n_1541 & ~n_1542;
assign n_1544 =  x_2117 & ~n_1513;
assign n_1545 =  i_27 &  n_1513;
assign n_1546 = ~n_1544 & ~n_1545;
assign n_1547 =  x_2117 & ~n_1546;
assign n_1548 = ~x_2117 &  n_1546;
assign n_1549 = ~n_1547 & ~n_1548;
assign n_1550 =  x_2116 & ~n_1513;
assign n_1551 =  i_26 &  n_1513;
assign n_1552 = ~n_1550 & ~n_1551;
assign n_1553 =  x_2116 & ~n_1552;
assign n_1554 = ~x_2116 &  n_1552;
assign n_1555 = ~n_1553 & ~n_1554;
assign n_1556 =  x_2115 & ~n_1513;
assign n_1557 =  i_25 &  n_1513;
assign n_1558 = ~n_1556 & ~n_1557;
assign n_1559 =  x_2115 & ~n_1558;
assign n_1560 = ~x_2115 &  n_1558;
assign n_1561 = ~n_1559 & ~n_1560;
assign n_1562 =  x_2114 & ~n_1513;
assign n_1563 =  i_24 &  n_1513;
assign n_1564 = ~n_1562 & ~n_1563;
assign n_1565 =  x_2114 & ~n_1564;
assign n_1566 = ~x_2114 &  n_1564;
assign n_1567 = ~n_1565 & ~n_1566;
assign n_1568 =  x_2113 & ~n_1513;
assign n_1569 =  i_23 &  n_1513;
assign n_1570 = ~n_1568 & ~n_1569;
assign n_1571 =  x_2113 & ~n_1570;
assign n_1572 = ~x_2113 &  n_1570;
assign n_1573 = ~n_1571 & ~n_1572;
assign n_1574 =  x_2112 & ~n_1513;
assign n_1575 =  i_22 &  n_1513;
assign n_1576 = ~n_1574 & ~n_1575;
assign n_1577 =  x_2112 & ~n_1576;
assign n_1578 = ~x_2112 &  n_1576;
assign n_1579 = ~n_1577 & ~n_1578;
assign n_1580 =  x_2111 & ~n_1513;
assign n_1581 =  i_21 &  n_1513;
assign n_1582 = ~n_1580 & ~n_1581;
assign n_1583 =  x_2111 & ~n_1582;
assign n_1584 = ~x_2111 &  n_1582;
assign n_1585 = ~n_1583 & ~n_1584;
assign n_1586 =  x_2110 & ~n_1513;
assign n_1587 =  i_20 &  n_1513;
assign n_1588 = ~n_1586 & ~n_1587;
assign n_1589 =  x_2110 & ~n_1588;
assign n_1590 = ~x_2110 &  n_1588;
assign n_1591 = ~n_1589 & ~n_1590;
assign n_1592 =  x_2109 & ~n_1513;
assign n_1593 =  i_19 &  n_1513;
assign n_1594 = ~n_1592 & ~n_1593;
assign n_1595 =  x_2109 & ~n_1594;
assign n_1596 = ~x_2109 &  n_1594;
assign n_1597 = ~n_1595 & ~n_1596;
assign n_1598 =  x_2108 & ~n_1513;
assign n_1599 =  i_18 &  n_1513;
assign n_1600 = ~n_1598 & ~n_1599;
assign n_1601 =  x_2108 & ~n_1600;
assign n_1602 = ~x_2108 &  n_1600;
assign n_1603 = ~n_1601 & ~n_1602;
assign n_1604 =  x_2107 & ~n_1513;
assign n_1605 =  i_17 &  n_1513;
assign n_1606 = ~n_1604 & ~n_1605;
assign n_1607 =  x_2107 & ~n_1606;
assign n_1608 = ~x_2107 &  n_1606;
assign n_1609 = ~n_1607 & ~n_1608;
assign n_1610 =  x_2106 & ~n_1513;
assign n_1611 =  i_16 &  n_1513;
assign n_1612 = ~n_1610 & ~n_1611;
assign n_1613 =  x_2106 & ~n_1612;
assign n_1614 = ~x_2106 &  n_1612;
assign n_1615 = ~n_1613 & ~n_1614;
assign n_1616 =  x_2105 & ~n_1513;
assign n_1617 =  i_15 &  n_1513;
assign n_1618 = ~n_1616 & ~n_1617;
assign n_1619 =  x_2105 & ~n_1618;
assign n_1620 = ~x_2105 &  n_1618;
assign n_1621 = ~n_1619 & ~n_1620;
assign n_1622 =  x_2104 & ~n_1513;
assign n_1623 =  i_14 &  n_1513;
assign n_1624 = ~n_1622 & ~n_1623;
assign n_1625 =  x_2104 & ~n_1624;
assign n_1626 = ~x_2104 &  n_1624;
assign n_1627 = ~n_1625 & ~n_1626;
assign n_1628 =  x_2103 & ~n_1513;
assign n_1629 =  i_13 &  n_1513;
assign n_1630 = ~n_1628 & ~n_1629;
assign n_1631 =  x_2103 & ~n_1630;
assign n_1632 = ~x_2103 &  n_1630;
assign n_1633 = ~n_1631 & ~n_1632;
assign n_1634 =  x_2102 & ~n_1513;
assign n_1635 =  i_12 &  n_1513;
assign n_1636 = ~n_1634 & ~n_1635;
assign n_1637 =  x_2102 & ~n_1636;
assign n_1638 = ~x_2102 &  n_1636;
assign n_1639 = ~n_1637 & ~n_1638;
assign n_1640 =  x_2101 & ~n_1513;
assign n_1641 =  i_11 &  n_1513;
assign n_1642 = ~n_1640 & ~n_1641;
assign n_1643 =  x_2101 & ~n_1642;
assign n_1644 = ~x_2101 &  n_1642;
assign n_1645 = ~n_1643 & ~n_1644;
assign n_1646 =  x_2100 & ~n_1513;
assign n_1647 =  i_10 &  n_1513;
assign n_1648 = ~n_1646 & ~n_1647;
assign n_1649 =  x_2100 & ~n_1648;
assign n_1650 = ~x_2100 &  n_1648;
assign n_1651 = ~n_1649 & ~n_1650;
assign n_1652 =  x_2099 & ~n_1513;
assign n_1653 =  i_9 &  n_1513;
assign n_1654 = ~n_1652 & ~n_1653;
assign n_1655 =  x_2099 & ~n_1654;
assign n_1656 = ~x_2099 &  n_1654;
assign n_1657 = ~n_1655 & ~n_1656;
assign n_1658 =  x_2098 & ~n_1513;
assign n_1659 =  i_8 &  n_1513;
assign n_1660 = ~n_1658 & ~n_1659;
assign n_1661 =  x_2098 & ~n_1660;
assign n_1662 = ~x_2098 &  n_1660;
assign n_1663 = ~n_1661 & ~n_1662;
assign n_1664 =  x_2097 & ~n_1513;
assign n_1665 =  i_7 &  n_1513;
assign n_1666 = ~n_1664 & ~n_1665;
assign n_1667 =  x_2097 & ~n_1666;
assign n_1668 = ~x_2097 &  n_1666;
assign n_1669 = ~n_1667 & ~n_1668;
assign n_1670 =  x_2096 & ~n_1513;
assign n_1671 =  i_6 &  n_1513;
assign n_1672 = ~n_1670 & ~n_1671;
assign n_1673 =  x_2096 & ~n_1672;
assign n_1674 = ~x_2096 &  n_1672;
assign n_1675 = ~n_1673 & ~n_1674;
assign n_1676 =  x_2095 & ~n_1513;
assign n_1677 =  i_5 &  n_1513;
assign n_1678 = ~n_1676 & ~n_1677;
assign n_1679 =  x_2095 & ~n_1678;
assign n_1680 = ~x_2095 &  n_1678;
assign n_1681 = ~n_1679 & ~n_1680;
assign n_1682 =  x_2094 & ~n_1513;
assign n_1683 =  i_4 &  n_1513;
assign n_1684 = ~n_1682 & ~n_1683;
assign n_1685 =  x_2094 & ~n_1684;
assign n_1686 = ~x_2094 &  n_1684;
assign n_1687 = ~n_1685 & ~n_1686;
assign n_1688 =  x_2093 & ~n_1513;
assign n_1689 =  i_3 &  n_1513;
assign n_1690 = ~n_1688 & ~n_1689;
assign n_1691 =  x_2093 & ~n_1690;
assign n_1692 = ~x_2093 &  n_1690;
assign n_1693 = ~n_1691 & ~n_1692;
assign n_1694 =  x_2092 & ~n_1513;
assign n_1695 =  i_2 &  n_1513;
assign n_1696 = ~n_1694 & ~n_1695;
assign n_1697 =  x_2092 & ~n_1696;
assign n_1698 = ~x_2092 &  n_1696;
assign n_1699 = ~n_1697 & ~n_1698;
assign n_1700 =  x_2091 & ~n_1513;
assign n_1701 =  i_1 &  n_1513;
assign n_1702 = ~n_1700 & ~n_1701;
assign n_1703 =  x_2091 & ~n_1702;
assign n_1704 = ~x_2091 &  n_1702;
assign n_1705 = ~n_1703 & ~n_1704;
assign n_1706 = ~x_41 & ~x_42;
assign n_1707 =  n_184 &  n_1706;
assign n_1708 = ~x_36 &  n_387;
assign n_1709 =  n_187 &  n_1708;
assign n_1710 =  n_1707 &  n_1709;
assign n_1711 =  x_2090 & ~n_1710;
assign n_1712 =  i_32 &  n_1710;
assign n_1713 = ~n_1711 & ~n_1712;
assign n_1714 =  x_2090 & ~n_1713;
assign n_1715 = ~x_2090 &  n_1713;
assign n_1716 = ~n_1714 & ~n_1715;
assign n_1717 =  x_2089 & ~n_1710;
assign n_1718 =  i_31 &  n_1710;
assign n_1719 = ~n_1717 & ~n_1718;
assign n_1720 =  x_2089 & ~n_1719;
assign n_1721 = ~x_2089 &  n_1719;
assign n_1722 = ~n_1720 & ~n_1721;
assign n_1723 =  x_2088 & ~n_1710;
assign n_1724 =  i_30 &  n_1710;
assign n_1725 = ~n_1723 & ~n_1724;
assign n_1726 =  x_2088 & ~n_1725;
assign n_1727 = ~x_2088 &  n_1725;
assign n_1728 = ~n_1726 & ~n_1727;
assign n_1729 =  x_2087 & ~n_1710;
assign n_1730 =  i_29 &  n_1710;
assign n_1731 = ~n_1729 & ~n_1730;
assign n_1732 =  x_2087 & ~n_1731;
assign n_1733 = ~x_2087 &  n_1731;
assign n_1734 = ~n_1732 & ~n_1733;
assign n_1735 =  x_2086 & ~n_1710;
assign n_1736 =  i_28 &  n_1710;
assign n_1737 = ~n_1735 & ~n_1736;
assign n_1738 =  x_2086 & ~n_1737;
assign n_1739 = ~x_2086 &  n_1737;
assign n_1740 = ~n_1738 & ~n_1739;
assign n_1741 =  x_2085 & ~n_1710;
assign n_1742 =  i_27 &  n_1710;
assign n_1743 = ~n_1741 & ~n_1742;
assign n_1744 =  x_2085 & ~n_1743;
assign n_1745 = ~x_2085 &  n_1743;
assign n_1746 = ~n_1744 & ~n_1745;
assign n_1747 =  x_2084 & ~n_1710;
assign n_1748 =  i_26 &  n_1710;
assign n_1749 = ~n_1747 & ~n_1748;
assign n_1750 =  x_2084 & ~n_1749;
assign n_1751 = ~x_2084 &  n_1749;
assign n_1752 = ~n_1750 & ~n_1751;
assign n_1753 =  x_2083 & ~n_1710;
assign n_1754 =  i_25 &  n_1710;
assign n_1755 = ~n_1753 & ~n_1754;
assign n_1756 =  x_2083 & ~n_1755;
assign n_1757 = ~x_2083 &  n_1755;
assign n_1758 = ~n_1756 & ~n_1757;
assign n_1759 =  x_2082 & ~n_1710;
assign n_1760 =  i_24 &  n_1710;
assign n_1761 = ~n_1759 & ~n_1760;
assign n_1762 =  x_2082 & ~n_1761;
assign n_1763 = ~x_2082 &  n_1761;
assign n_1764 = ~n_1762 & ~n_1763;
assign n_1765 =  x_2081 & ~n_1710;
assign n_1766 =  i_23 &  n_1710;
assign n_1767 = ~n_1765 & ~n_1766;
assign n_1768 =  x_2081 & ~n_1767;
assign n_1769 = ~x_2081 &  n_1767;
assign n_1770 = ~n_1768 & ~n_1769;
assign n_1771 =  x_2080 & ~n_1710;
assign n_1772 =  i_22 &  n_1710;
assign n_1773 = ~n_1771 & ~n_1772;
assign n_1774 =  x_2080 & ~n_1773;
assign n_1775 = ~x_2080 &  n_1773;
assign n_1776 = ~n_1774 & ~n_1775;
assign n_1777 =  x_2079 & ~n_1710;
assign n_1778 =  i_21 &  n_1710;
assign n_1779 = ~n_1777 & ~n_1778;
assign n_1780 =  x_2079 & ~n_1779;
assign n_1781 = ~x_2079 &  n_1779;
assign n_1782 = ~n_1780 & ~n_1781;
assign n_1783 =  x_2078 & ~n_1710;
assign n_1784 =  i_20 &  n_1710;
assign n_1785 = ~n_1783 & ~n_1784;
assign n_1786 =  x_2078 & ~n_1785;
assign n_1787 = ~x_2078 &  n_1785;
assign n_1788 = ~n_1786 & ~n_1787;
assign n_1789 =  x_2077 & ~n_1710;
assign n_1790 =  i_19 &  n_1710;
assign n_1791 = ~n_1789 & ~n_1790;
assign n_1792 =  x_2077 & ~n_1791;
assign n_1793 = ~x_2077 &  n_1791;
assign n_1794 = ~n_1792 & ~n_1793;
assign n_1795 =  x_2076 & ~n_1710;
assign n_1796 =  i_18 &  n_1710;
assign n_1797 = ~n_1795 & ~n_1796;
assign n_1798 =  x_2076 & ~n_1797;
assign n_1799 = ~x_2076 &  n_1797;
assign n_1800 = ~n_1798 & ~n_1799;
assign n_1801 =  x_2075 & ~n_1710;
assign n_1802 =  i_17 &  n_1710;
assign n_1803 = ~n_1801 & ~n_1802;
assign n_1804 =  x_2075 & ~n_1803;
assign n_1805 = ~x_2075 &  n_1803;
assign n_1806 = ~n_1804 & ~n_1805;
assign n_1807 =  x_2074 & ~n_1710;
assign n_1808 =  i_16 &  n_1710;
assign n_1809 = ~n_1807 & ~n_1808;
assign n_1810 =  x_2074 & ~n_1809;
assign n_1811 = ~x_2074 &  n_1809;
assign n_1812 = ~n_1810 & ~n_1811;
assign n_1813 =  x_2073 & ~n_1710;
assign n_1814 =  i_15 &  n_1710;
assign n_1815 = ~n_1813 & ~n_1814;
assign n_1816 =  x_2073 & ~n_1815;
assign n_1817 = ~x_2073 &  n_1815;
assign n_1818 = ~n_1816 & ~n_1817;
assign n_1819 =  x_2072 & ~n_1710;
assign n_1820 =  i_14 &  n_1710;
assign n_1821 = ~n_1819 & ~n_1820;
assign n_1822 =  x_2072 & ~n_1821;
assign n_1823 = ~x_2072 &  n_1821;
assign n_1824 = ~n_1822 & ~n_1823;
assign n_1825 =  x_2071 & ~n_1710;
assign n_1826 =  i_13 &  n_1710;
assign n_1827 = ~n_1825 & ~n_1826;
assign n_1828 =  x_2071 & ~n_1827;
assign n_1829 = ~x_2071 &  n_1827;
assign n_1830 = ~n_1828 & ~n_1829;
assign n_1831 =  x_2070 & ~n_1710;
assign n_1832 =  i_12 &  n_1710;
assign n_1833 = ~n_1831 & ~n_1832;
assign n_1834 =  x_2070 & ~n_1833;
assign n_1835 = ~x_2070 &  n_1833;
assign n_1836 = ~n_1834 & ~n_1835;
assign n_1837 =  x_2069 & ~n_1710;
assign n_1838 =  i_11 &  n_1710;
assign n_1839 = ~n_1837 & ~n_1838;
assign n_1840 =  x_2069 & ~n_1839;
assign n_1841 = ~x_2069 &  n_1839;
assign n_1842 = ~n_1840 & ~n_1841;
assign n_1843 =  x_2068 & ~n_1710;
assign n_1844 =  i_10 &  n_1710;
assign n_1845 = ~n_1843 & ~n_1844;
assign n_1846 =  x_2068 & ~n_1845;
assign n_1847 = ~x_2068 &  n_1845;
assign n_1848 = ~n_1846 & ~n_1847;
assign n_1849 =  x_2067 & ~n_1710;
assign n_1850 =  i_9 &  n_1710;
assign n_1851 = ~n_1849 & ~n_1850;
assign n_1852 =  x_2067 & ~n_1851;
assign n_1853 = ~x_2067 &  n_1851;
assign n_1854 = ~n_1852 & ~n_1853;
assign n_1855 =  x_2066 & ~n_1710;
assign n_1856 =  i_8 &  n_1710;
assign n_1857 = ~n_1855 & ~n_1856;
assign n_1858 =  x_2066 & ~n_1857;
assign n_1859 = ~x_2066 &  n_1857;
assign n_1860 = ~n_1858 & ~n_1859;
assign n_1861 =  x_2065 & ~n_1710;
assign n_1862 =  i_7 &  n_1710;
assign n_1863 = ~n_1861 & ~n_1862;
assign n_1864 =  x_2065 & ~n_1863;
assign n_1865 = ~x_2065 &  n_1863;
assign n_1866 = ~n_1864 & ~n_1865;
assign n_1867 =  x_2064 & ~n_1710;
assign n_1868 =  i_6 &  n_1710;
assign n_1869 = ~n_1867 & ~n_1868;
assign n_1870 =  x_2064 & ~n_1869;
assign n_1871 = ~x_2064 &  n_1869;
assign n_1872 = ~n_1870 & ~n_1871;
assign n_1873 =  x_2063 & ~n_1710;
assign n_1874 =  i_5 &  n_1710;
assign n_1875 = ~n_1873 & ~n_1874;
assign n_1876 =  x_2063 & ~n_1875;
assign n_1877 = ~x_2063 &  n_1875;
assign n_1878 = ~n_1876 & ~n_1877;
assign n_1879 =  x_2062 & ~n_1710;
assign n_1880 =  i_4 &  n_1710;
assign n_1881 = ~n_1879 & ~n_1880;
assign n_1882 =  x_2062 & ~n_1881;
assign n_1883 = ~x_2062 &  n_1881;
assign n_1884 = ~n_1882 & ~n_1883;
assign n_1885 =  x_2061 & ~n_1710;
assign n_1886 =  i_3 &  n_1710;
assign n_1887 = ~n_1885 & ~n_1886;
assign n_1888 =  x_2061 & ~n_1887;
assign n_1889 = ~x_2061 &  n_1887;
assign n_1890 = ~n_1888 & ~n_1889;
assign n_1891 =  x_2060 & ~n_1710;
assign n_1892 =  i_2 &  n_1710;
assign n_1893 = ~n_1891 & ~n_1892;
assign n_1894 =  x_2060 & ~n_1893;
assign n_1895 = ~x_2060 &  n_1893;
assign n_1896 = ~n_1894 & ~n_1895;
assign n_1897 =  x_2059 & ~n_1710;
assign n_1898 =  i_1 &  n_1710;
assign n_1899 = ~n_1897 & ~n_1898;
assign n_1900 =  x_2059 & ~n_1899;
assign n_1901 = ~x_2059 &  n_1899;
assign n_1902 = ~n_1900 & ~n_1901;
assign n_1903 = ~x_36 &  n_981;
assign n_1904 =  n_389 &  n_1903;
assign n_1905 = ~x_39 &  n_585;
assign n_1906 = ~x_42 &  n_1905;
assign n_1907 =  n_1904 &  n_1906;
assign n_1908 =  x_2058 & ~n_1907;
assign n_1909 =  i_32 &  n_1907;
assign n_1910 = ~n_1908 & ~n_1909;
assign n_1911 =  x_2058 & ~n_1910;
assign n_1912 = ~x_2058 &  n_1910;
assign n_1913 = ~n_1911 & ~n_1912;
assign n_1914 =  x_2057 & ~n_1907;
assign n_1915 =  i_31 &  n_1907;
assign n_1916 = ~n_1914 & ~n_1915;
assign n_1917 =  x_2057 & ~n_1916;
assign n_1918 = ~x_2057 &  n_1916;
assign n_1919 = ~n_1917 & ~n_1918;
assign n_1920 =  x_2056 & ~n_1907;
assign n_1921 =  i_30 &  n_1907;
assign n_1922 = ~n_1920 & ~n_1921;
assign n_1923 =  x_2056 & ~n_1922;
assign n_1924 = ~x_2056 &  n_1922;
assign n_1925 = ~n_1923 & ~n_1924;
assign n_1926 =  x_2055 & ~n_1907;
assign n_1927 =  i_29 &  n_1907;
assign n_1928 = ~n_1926 & ~n_1927;
assign n_1929 =  x_2055 & ~n_1928;
assign n_1930 = ~x_2055 &  n_1928;
assign n_1931 = ~n_1929 & ~n_1930;
assign n_1932 =  x_2054 & ~n_1907;
assign n_1933 =  i_28 &  n_1907;
assign n_1934 = ~n_1932 & ~n_1933;
assign n_1935 =  x_2054 & ~n_1934;
assign n_1936 = ~x_2054 &  n_1934;
assign n_1937 = ~n_1935 & ~n_1936;
assign n_1938 =  x_2053 & ~n_1907;
assign n_1939 =  i_27 &  n_1907;
assign n_1940 = ~n_1938 & ~n_1939;
assign n_1941 =  x_2053 & ~n_1940;
assign n_1942 = ~x_2053 &  n_1940;
assign n_1943 = ~n_1941 & ~n_1942;
assign n_1944 =  x_2052 & ~n_1907;
assign n_1945 =  i_26 &  n_1907;
assign n_1946 = ~n_1944 & ~n_1945;
assign n_1947 =  x_2052 & ~n_1946;
assign n_1948 = ~x_2052 &  n_1946;
assign n_1949 = ~n_1947 & ~n_1948;
assign n_1950 =  x_2051 & ~n_1907;
assign n_1951 =  i_25 &  n_1907;
assign n_1952 = ~n_1950 & ~n_1951;
assign n_1953 =  x_2051 & ~n_1952;
assign n_1954 = ~x_2051 &  n_1952;
assign n_1955 = ~n_1953 & ~n_1954;
assign n_1956 =  x_2050 & ~n_1907;
assign n_1957 =  i_24 &  n_1907;
assign n_1958 = ~n_1956 & ~n_1957;
assign n_1959 =  x_2050 & ~n_1958;
assign n_1960 = ~x_2050 &  n_1958;
assign n_1961 = ~n_1959 & ~n_1960;
assign n_1962 =  x_2049 & ~n_1907;
assign n_1963 =  i_23 &  n_1907;
assign n_1964 = ~n_1962 & ~n_1963;
assign n_1965 =  x_2049 & ~n_1964;
assign n_1966 = ~x_2049 &  n_1964;
assign n_1967 = ~n_1965 & ~n_1966;
assign n_1968 =  x_2048 & ~n_1907;
assign n_1969 =  i_22 &  n_1907;
assign n_1970 = ~n_1968 & ~n_1969;
assign n_1971 =  x_2048 & ~n_1970;
assign n_1972 = ~x_2048 &  n_1970;
assign n_1973 = ~n_1971 & ~n_1972;
assign n_1974 =  x_2047 & ~n_1907;
assign n_1975 =  i_21 &  n_1907;
assign n_1976 = ~n_1974 & ~n_1975;
assign n_1977 =  x_2047 & ~n_1976;
assign n_1978 = ~x_2047 &  n_1976;
assign n_1979 = ~n_1977 & ~n_1978;
assign n_1980 =  x_2046 & ~n_1907;
assign n_1981 =  i_20 &  n_1907;
assign n_1982 = ~n_1980 & ~n_1981;
assign n_1983 =  x_2046 & ~n_1982;
assign n_1984 = ~x_2046 &  n_1982;
assign n_1985 = ~n_1983 & ~n_1984;
assign n_1986 =  x_2045 & ~n_1907;
assign n_1987 =  i_19 &  n_1907;
assign n_1988 = ~n_1986 & ~n_1987;
assign n_1989 =  x_2045 & ~n_1988;
assign n_1990 = ~x_2045 &  n_1988;
assign n_1991 = ~n_1989 & ~n_1990;
assign n_1992 =  x_2044 & ~n_1907;
assign n_1993 =  i_18 &  n_1907;
assign n_1994 = ~n_1992 & ~n_1993;
assign n_1995 =  x_2044 & ~n_1994;
assign n_1996 = ~x_2044 &  n_1994;
assign n_1997 = ~n_1995 & ~n_1996;
assign n_1998 =  x_2043 & ~n_1907;
assign n_1999 =  i_17 &  n_1907;
assign n_2000 = ~n_1998 & ~n_1999;
assign n_2001 =  x_2043 & ~n_2000;
assign n_2002 = ~x_2043 &  n_2000;
assign n_2003 = ~n_2001 & ~n_2002;
assign n_2004 =  x_2042 & ~n_1907;
assign n_2005 =  i_16 &  n_1907;
assign n_2006 = ~n_2004 & ~n_2005;
assign n_2007 =  x_2042 & ~n_2006;
assign n_2008 = ~x_2042 &  n_2006;
assign n_2009 = ~n_2007 & ~n_2008;
assign n_2010 =  x_2041 & ~n_1907;
assign n_2011 =  i_15 &  n_1907;
assign n_2012 = ~n_2010 & ~n_2011;
assign n_2013 =  x_2041 & ~n_2012;
assign n_2014 = ~x_2041 &  n_2012;
assign n_2015 = ~n_2013 & ~n_2014;
assign n_2016 =  x_2040 & ~n_1907;
assign n_2017 =  i_14 &  n_1907;
assign n_2018 = ~n_2016 & ~n_2017;
assign n_2019 =  x_2040 & ~n_2018;
assign n_2020 = ~x_2040 &  n_2018;
assign n_2021 = ~n_2019 & ~n_2020;
assign n_2022 =  x_2039 & ~n_1907;
assign n_2023 =  i_13 &  n_1907;
assign n_2024 = ~n_2022 & ~n_2023;
assign n_2025 =  x_2039 & ~n_2024;
assign n_2026 = ~x_2039 &  n_2024;
assign n_2027 = ~n_2025 & ~n_2026;
assign n_2028 =  x_2038 & ~n_1907;
assign n_2029 =  i_12 &  n_1907;
assign n_2030 = ~n_2028 & ~n_2029;
assign n_2031 =  x_2038 & ~n_2030;
assign n_2032 = ~x_2038 &  n_2030;
assign n_2033 = ~n_2031 & ~n_2032;
assign n_2034 =  x_2037 & ~n_1907;
assign n_2035 =  i_11 &  n_1907;
assign n_2036 = ~n_2034 & ~n_2035;
assign n_2037 =  x_2037 & ~n_2036;
assign n_2038 = ~x_2037 &  n_2036;
assign n_2039 = ~n_2037 & ~n_2038;
assign n_2040 =  x_2036 & ~n_1907;
assign n_2041 =  i_10 &  n_1907;
assign n_2042 = ~n_2040 & ~n_2041;
assign n_2043 =  x_2036 & ~n_2042;
assign n_2044 = ~x_2036 &  n_2042;
assign n_2045 = ~n_2043 & ~n_2044;
assign n_2046 =  x_2035 & ~n_1907;
assign n_2047 =  i_9 &  n_1907;
assign n_2048 = ~n_2046 & ~n_2047;
assign n_2049 =  x_2035 & ~n_2048;
assign n_2050 = ~x_2035 &  n_2048;
assign n_2051 = ~n_2049 & ~n_2050;
assign n_2052 =  x_2034 & ~n_1907;
assign n_2053 =  i_8 &  n_1907;
assign n_2054 = ~n_2052 & ~n_2053;
assign n_2055 =  x_2034 & ~n_2054;
assign n_2056 = ~x_2034 &  n_2054;
assign n_2057 = ~n_2055 & ~n_2056;
assign n_2058 =  x_2033 & ~n_1907;
assign n_2059 =  i_7 &  n_1907;
assign n_2060 = ~n_2058 & ~n_2059;
assign n_2061 =  x_2033 & ~n_2060;
assign n_2062 = ~x_2033 &  n_2060;
assign n_2063 = ~n_2061 & ~n_2062;
assign n_2064 =  x_2032 & ~n_1907;
assign n_2065 =  i_6 &  n_1907;
assign n_2066 = ~n_2064 & ~n_2065;
assign n_2067 =  x_2032 & ~n_2066;
assign n_2068 = ~x_2032 &  n_2066;
assign n_2069 = ~n_2067 & ~n_2068;
assign n_2070 =  x_2031 & ~n_1907;
assign n_2071 =  i_5 &  n_1907;
assign n_2072 = ~n_2070 & ~n_2071;
assign n_2073 =  x_2031 & ~n_2072;
assign n_2074 = ~x_2031 &  n_2072;
assign n_2075 = ~n_2073 & ~n_2074;
assign n_2076 =  x_2030 & ~n_1907;
assign n_2077 =  i_4 &  n_1907;
assign n_2078 = ~n_2076 & ~n_2077;
assign n_2079 =  x_2030 & ~n_2078;
assign n_2080 = ~x_2030 &  n_2078;
assign n_2081 = ~n_2079 & ~n_2080;
assign n_2082 =  x_2029 & ~n_1907;
assign n_2083 =  i_3 &  n_1907;
assign n_2084 = ~n_2082 & ~n_2083;
assign n_2085 =  x_2029 & ~n_2084;
assign n_2086 = ~x_2029 &  n_2084;
assign n_2087 = ~n_2085 & ~n_2086;
assign n_2088 =  x_2028 & ~n_1907;
assign n_2089 =  i_2 &  n_1907;
assign n_2090 = ~n_2088 & ~n_2089;
assign n_2091 =  x_2028 & ~n_2090;
assign n_2092 = ~x_2028 &  n_2090;
assign n_2093 = ~n_2091 & ~n_2092;
assign n_2094 =  x_2027 & ~n_1907;
assign n_2095 =  i_1 &  n_1907;
assign n_2096 = ~n_2094 & ~n_2095;
assign n_2097 =  x_2027 & ~n_2096;
assign n_2098 = ~x_2027 &  n_2096;
assign n_2099 = ~n_2097 & ~n_2098;
assign n_2100 = ~x_37 & ~x_38;
assign n_2101 =  n_2100 &  n_190;
assign n_2102 =  n_186 &  n_2101;
assign n_2103 =  x_2026 & ~n_2102;
assign n_2104 =  i_32 &  n_2102;
assign n_2105 = ~n_2103 & ~n_2104;
assign n_2106 =  x_2026 & ~n_2105;
assign n_2107 = ~x_2026 &  n_2105;
assign n_2108 = ~n_2106 & ~n_2107;
assign n_2109 =  x_2025 & ~n_2102;
assign n_2110 =  i_31 &  n_2102;
assign n_2111 = ~n_2109 & ~n_2110;
assign n_2112 =  x_2025 & ~n_2111;
assign n_2113 = ~x_2025 &  n_2111;
assign n_2114 = ~n_2112 & ~n_2113;
assign n_2115 =  x_2024 & ~n_2102;
assign n_2116 =  i_30 &  n_2102;
assign n_2117 = ~n_2115 & ~n_2116;
assign n_2118 =  x_2024 & ~n_2117;
assign n_2119 = ~x_2024 &  n_2117;
assign n_2120 = ~n_2118 & ~n_2119;
assign n_2121 =  x_2023 & ~n_2102;
assign n_2122 =  i_29 &  n_2102;
assign n_2123 = ~n_2121 & ~n_2122;
assign n_2124 =  x_2023 & ~n_2123;
assign n_2125 = ~x_2023 &  n_2123;
assign n_2126 = ~n_2124 & ~n_2125;
assign n_2127 =  x_2022 & ~n_2102;
assign n_2128 =  i_28 &  n_2102;
assign n_2129 = ~n_2127 & ~n_2128;
assign n_2130 =  x_2022 & ~n_2129;
assign n_2131 = ~x_2022 &  n_2129;
assign n_2132 = ~n_2130 & ~n_2131;
assign n_2133 =  x_2021 & ~n_2102;
assign n_2134 =  i_27 &  n_2102;
assign n_2135 = ~n_2133 & ~n_2134;
assign n_2136 =  x_2021 & ~n_2135;
assign n_2137 = ~x_2021 &  n_2135;
assign n_2138 = ~n_2136 & ~n_2137;
assign n_2139 =  x_2020 & ~n_2102;
assign n_2140 =  i_26 &  n_2102;
assign n_2141 = ~n_2139 & ~n_2140;
assign n_2142 =  x_2020 & ~n_2141;
assign n_2143 = ~x_2020 &  n_2141;
assign n_2144 = ~n_2142 & ~n_2143;
assign n_2145 =  x_2019 & ~n_2102;
assign n_2146 =  i_25 &  n_2102;
assign n_2147 = ~n_2145 & ~n_2146;
assign n_2148 =  x_2019 & ~n_2147;
assign n_2149 = ~x_2019 &  n_2147;
assign n_2150 = ~n_2148 & ~n_2149;
assign n_2151 =  x_2018 & ~n_2102;
assign n_2152 =  i_24 &  n_2102;
assign n_2153 = ~n_2151 & ~n_2152;
assign n_2154 =  x_2018 & ~n_2153;
assign n_2155 = ~x_2018 &  n_2153;
assign n_2156 = ~n_2154 & ~n_2155;
assign n_2157 =  x_2017 & ~n_2102;
assign n_2158 =  i_23 &  n_2102;
assign n_2159 = ~n_2157 & ~n_2158;
assign n_2160 =  x_2017 & ~n_2159;
assign n_2161 = ~x_2017 &  n_2159;
assign n_2162 = ~n_2160 & ~n_2161;
assign n_2163 =  x_2016 & ~n_2102;
assign n_2164 =  i_22 &  n_2102;
assign n_2165 = ~n_2163 & ~n_2164;
assign n_2166 =  x_2016 & ~n_2165;
assign n_2167 = ~x_2016 &  n_2165;
assign n_2168 = ~n_2166 & ~n_2167;
assign n_2169 =  x_2015 & ~n_2102;
assign n_2170 =  i_21 &  n_2102;
assign n_2171 = ~n_2169 & ~n_2170;
assign n_2172 =  x_2015 & ~n_2171;
assign n_2173 = ~x_2015 &  n_2171;
assign n_2174 = ~n_2172 & ~n_2173;
assign n_2175 =  x_2014 & ~n_2102;
assign n_2176 =  i_20 &  n_2102;
assign n_2177 = ~n_2175 & ~n_2176;
assign n_2178 =  x_2014 & ~n_2177;
assign n_2179 = ~x_2014 &  n_2177;
assign n_2180 = ~n_2178 & ~n_2179;
assign n_2181 =  x_2013 & ~n_2102;
assign n_2182 =  i_19 &  n_2102;
assign n_2183 = ~n_2181 & ~n_2182;
assign n_2184 =  x_2013 & ~n_2183;
assign n_2185 = ~x_2013 &  n_2183;
assign n_2186 = ~n_2184 & ~n_2185;
assign n_2187 =  x_2012 & ~n_2102;
assign n_2188 =  i_18 &  n_2102;
assign n_2189 = ~n_2187 & ~n_2188;
assign n_2190 =  x_2012 & ~n_2189;
assign n_2191 = ~x_2012 &  n_2189;
assign n_2192 = ~n_2190 & ~n_2191;
assign n_2193 =  x_2011 & ~n_2102;
assign n_2194 =  i_17 &  n_2102;
assign n_2195 = ~n_2193 & ~n_2194;
assign n_2196 =  x_2011 & ~n_2195;
assign n_2197 = ~x_2011 &  n_2195;
assign n_2198 = ~n_2196 & ~n_2197;
assign n_2199 =  x_2010 & ~n_2102;
assign n_2200 =  i_16 &  n_2102;
assign n_2201 = ~n_2199 & ~n_2200;
assign n_2202 =  x_2010 & ~n_2201;
assign n_2203 = ~x_2010 &  n_2201;
assign n_2204 = ~n_2202 & ~n_2203;
assign n_2205 =  x_2009 & ~n_2102;
assign n_2206 =  i_15 &  n_2102;
assign n_2207 = ~n_2205 & ~n_2206;
assign n_2208 =  x_2009 & ~n_2207;
assign n_2209 = ~x_2009 &  n_2207;
assign n_2210 = ~n_2208 & ~n_2209;
assign n_2211 =  x_2008 & ~n_2102;
assign n_2212 =  i_14 &  n_2102;
assign n_2213 = ~n_2211 & ~n_2212;
assign n_2214 =  x_2008 & ~n_2213;
assign n_2215 = ~x_2008 &  n_2213;
assign n_2216 = ~n_2214 & ~n_2215;
assign n_2217 =  x_2007 & ~n_2102;
assign n_2218 =  i_13 &  n_2102;
assign n_2219 = ~n_2217 & ~n_2218;
assign n_2220 =  x_2007 & ~n_2219;
assign n_2221 = ~x_2007 &  n_2219;
assign n_2222 = ~n_2220 & ~n_2221;
assign n_2223 =  x_2006 & ~n_2102;
assign n_2224 =  i_12 &  n_2102;
assign n_2225 = ~n_2223 & ~n_2224;
assign n_2226 =  x_2006 & ~n_2225;
assign n_2227 = ~x_2006 &  n_2225;
assign n_2228 = ~n_2226 & ~n_2227;
assign n_2229 =  x_2005 & ~n_2102;
assign n_2230 =  i_11 &  n_2102;
assign n_2231 = ~n_2229 & ~n_2230;
assign n_2232 =  x_2005 & ~n_2231;
assign n_2233 = ~x_2005 &  n_2231;
assign n_2234 = ~n_2232 & ~n_2233;
assign n_2235 =  x_2004 & ~n_2102;
assign n_2236 =  i_10 &  n_2102;
assign n_2237 = ~n_2235 & ~n_2236;
assign n_2238 =  x_2004 & ~n_2237;
assign n_2239 = ~x_2004 &  n_2237;
assign n_2240 = ~n_2238 & ~n_2239;
assign n_2241 =  x_2003 & ~n_2102;
assign n_2242 =  i_9 &  n_2102;
assign n_2243 = ~n_2241 & ~n_2242;
assign n_2244 =  x_2003 & ~n_2243;
assign n_2245 = ~x_2003 &  n_2243;
assign n_2246 = ~n_2244 & ~n_2245;
assign n_2247 =  x_2002 & ~n_2102;
assign n_2248 =  i_8 &  n_2102;
assign n_2249 = ~n_2247 & ~n_2248;
assign n_2250 =  x_2002 & ~n_2249;
assign n_2251 = ~x_2002 &  n_2249;
assign n_2252 = ~n_2250 & ~n_2251;
assign n_2253 =  x_2001 & ~n_2102;
assign n_2254 =  i_7 &  n_2102;
assign n_2255 = ~n_2253 & ~n_2254;
assign n_2256 =  x_2001 & ~n_2255;
assign n_2257 = ~x_2001 &  n_2255;
assign n_2258 = ~n_2256 & ~n_2257;
assign n_2259 =  x_2000 & ~n_2102;
assign n_2260 =  i_6 &  n_2102;
assign n_2261 = ~n_2259 & ~n_2260;
assign n_2262 =  x_2000 & ~n_2261;
assign n_2263 = ~x_2000 &  n_2261;
assign n_2264 = ~n_2262 & ~n_2263;
assign n_2265 =  x_1999 & ~n_2102;
assign n_2266 =  i_5 &  n_2102;
assign n_2267 = ~n_2265 & ~n_2266;
assign n_2268 =  x_1999 & ~n_2267;
assign n_2269 = ~x_1999 &  n_2267;
assign n_2270 = ~n_2268 & ~n_2269;
assign n_2271 =  x_1998 & ~n_2102;
assign n_2272 =  i_4 &  n_2102;
assign n_2273 = ~n_2271 & ~n_2272;
assign n_2274 =  x_1998 & ~n_2273;
assign n_2275 = ~x_1998 &  n_2273;
assign n_2276 = ~n_2274 & ~n_2275;
assign n_2277 =  x_1997 & ~n_2102;
assign n_2278 =  i_3 &  n_2102;
assign n_2279 = ~n_2277 & ~n_2278;
assign n_2280 =  x_1997 & ~n_2279;
assign n_2281 = ~x_1997 &  n_2279;
assign n_2282 = ~n_2280 & ~n_2281;
assign n_2283 =  x_1996 & ~n_2102;
assign n_2284 =  i_2 &  n_2102;
assign n_2285 = ~n_2283 & ~n_2284;
assign n_2286 =  x_1996 & ~n_2285;
assign n_2287 = ~x_1996 &  n_2285;
assign n_2288 = ~n_2286 & ~n_2287;
assign n_2289 =  x_1995 & ~n_2102;
assign n_2290 =  i_1 &  n_2102;
assign n_2291 = ~n_2289 & ~n_2290;
assign n_2292 =  x_1995 & ~n_2291;
assign n_2293 = ~x_1995 &  n_2291;
assign n_2294 = ~n_2292 & ~n_2293;
assign n_2295 = ~x_36 & ~x_37;
assign n_2296 =  n_2295 &  n_387;
assign n_2297 = ~x_38 &  n_2296;
assign n_2298 =  x_39 &  x_40;
assign n_2299 = ~x_41 &  n_2298;
assign n_2300 =  n_2297 &  n_2299;
assign n_2301 =  x_40 &  x_41;
assign n_2302 = ~x_39 &  n_187;
assign n_2303 =  n_982 &  n_2302;
assign n_2304 =  n_2301 &  n_2303;
assign n_2305 = ~n_2300 & ~n_2304;
assign n_2306 =  x_42 & ~n_2305;
assign n_2307 =  x_1994 & ~n_2306;
assign n_2308 =  i_32 &  n_2306;
assign n_2309 = ~n_2307 & ~n_2308;
assign n_2310 =  x_1994 & ~n_2309;
assign n_2311 = ~x_1994 &  n_2309;
assign n_2312 = ~n_2310 & ~n_2311;
assign n_2313 =  x_1993 & ~n_2306;
assign n_2314 =  i_31 &  n_2306;
assign n_2315 = ~n_2313 & ~n_2314;
assign n_2316 =  x_1993 & ~n_2315;
assign n_2317 = ~x_1993 &  n_2315;
assign n_2318 = ~n_2316 & ~n_2317;
assign n_2319 =  x_1992 & ~n_2306;
assign n_2320 =  i_30 &  n_2306;
assign n_2321 = ~n_2319 & ~n_2320;
assign n_2322 =  x_1992 & ~n_2321;
assign n_2323 = ~x_1992 &  n_2321;
assign n_2324 = ~n_2322 & ~n_2323;
assign n_2325 =  x_1991 & ~n_2306;
assign n_2326 =  i_29 &  n_2306;
assign n_2327 = ~n_2325 & ~n_2326;
assign n_2328 =  x_1991 & ~n_2327;
assign n_2329 = ~x_1991 &  n_2327;
assign n_2330 = ~n_2328 & ~n_2329;
assign n_2331 =  x_1990 & ~n_2306;
assign n_2332 =  i_28 &  n_2306;
assign n_2333 = ~n_2331 & ~n_2332;
assign n_2334 =  x_1990 & ~n_2333;
assign n_2335 = ~x_1990 &  n_2333;
assign n_2336 = ~n_2334 & ~n_2335;
assign n_2337 =  x_1989 & ~n_2306;
assign n_2338 =  i_27 &  n_2306;
assign n_2339 = ~n_2337 & ~n_2338;
assign n_2340 =  x_1989 & ~n_2339;
assign n_2341 = ~x_1989 &  n_2339;
assign n_2342 = ~n_2340 & ~n_2341;
assign n_2343 =  x_1988 & ~n_2306;
assign n_2344 =  i_26 &  n_2306;
assign n_2345 = ~n_2343 & ~n_2344;
assign n_2346 =  x_1988 & ~n_2345;
assign n_2347 = ~x_1988 &  n_2345;
assign n_2348 = ~n_2346 & ~n_2347;
assign n_2349 =  x_1987 & ~n_2306;
assign n_2350 =  i_25 &  n_2306;
assign n_2351 = ~n_2349 & ~n_2350;
assign n_2352 =  x_1987 & ~n_2351;
assign n_2353 = ~x_1987 &  n_2351;
assign n_2354 = ~n_2352 & ~n_2353;
assign n_2355 =  x_1986 & ~n_2306;
assign n_2356 =  i_24 &  n_2306;
assign n_2357 = ~n_2355 & ~n_2356;
assign n_2358 =  x_1986 & ~n_2357;
assign n_2359 = ~x_1986 &  n_2357;
assign n_2360 = ~n_2358 & ~n_2359;
assign n_2361 =  x_1985 & ~n_2306;
assign n_2362 =  i_23 &  n_2306;
assign n_2363 = ~n_2361 & ~n_2362;
assign n_2364 =  x_1985 & ~n_2363;
assign n_2365 = ~x_1985 &  n_2363;
assign n_2366 = ~n_2364 & ~n_2365;
assign n_2367 =  x_1984 & ~n_2306;
assign n_2368 =  i_22 &  n_2306;
assign n_2369 = ~n_2367 & ~n_2368;
assign n_2370 =  x_1984 & ~n_2369;
assign n_2371 = ~x_1984 &  n_2369;
assign n_2372 = ~n_2370 & ~n_2371;
assign n_2373 =  x_1983 & ~n_2306;
assign n_2374 =  i_21 &  n_2306;
assign n_2375 = ~n_2373 & ~n_2374;
assign n_2376 =  x_1983 & ~n_2375;
assign n_2377 = ~x_1983 &  n_2375;
assign n_2378 = ~n_2376 & ~n_2377;
assign n_2379 =  x_1982 & ~n_2306;
assign n_2380 =  i_20 &  n_2306;
assign n_2381 = ~n_2379 & ~n_2380;
assign n_2382 =  x_1982 & ~n_2381;
assign n_2383 = ~x_1982 &  n_2381;
assign n_2384 = ~n_2382 & ~n_2383;
assign n_2385 =  x_1981 & ~n_2306;
assign n_2386 =  i_19 &  n_2306;
assign n_2387 = ~n_2385 & ~n_2386;
assign n_2388 =  x_1981 & ~n_2387;
assign n_2389 = ~x_1981 &  n_2387;
assign n_2390 = ~n_2388 & ~n_2389;
assign n_2391 =  x_1980 & ~n_2306;
assign n_2392 =  i_18 &  n_2306;
assign n_2393 = ~n_2391 & ~n_2392;
assign n_2394 =  x_1980 & ~n_2393;
assign n_2395 = ~x_1980 &  n_2393;
assign n_2396 = ~n_2394 & ~n_2395;
assign n_2397 =  x_1979 & ~n_2306;
assign n_2398 =  i_17 &  n_2306;
assign n_2399 = ~n_2397 & ~n_2398;
assign n_2400 =  x_1979 & ~n_2399;
assign n_2401 = ~x_1979 &  n_2399;
assign n_2402 = ~n_2400 & ~n_2401;
assign n_2403 =  x_1978 & ~n_2306;
assign n_2404 =  i_16 &  n_2306;
assign n_2405 = ~n_2403 & ~n_2404;
assign n_2406 =  x_1978 & ~n_2405;
assign n_2407 = ~x_1978 &  n_2405;
assign n_2408 = ~n_2406 & ~n_2407;
assign n_2409 =  x_1977 & ~n_2306;
assign n_2410 =  i_15 &  n_2306;
assign n_2411 = ~n_2409 & ~n_2410;
assign n_2412 =  x_1977 & ~n_2411;
assign n_2413 = ~x_1977 &  n_2411;
assign n_2414 = ~n_2412 & ~n_2413;
assign n_2415 =  x_1976 & ~n_2306;
assign n_2416 =  i_14 &  n_2306;
assign n_2417 = ~n_2415 & ~n_2416;
assign n_2418 =  x_1976 & ~n_2417;
assign n_2419 = ~x_1976 &  n_2417;
assign n_2420 = ~n_2418 & ~n_2419;
assign n_2421 =  x_1975 & ~n_2306;
assign n_2422 =  i_13 &  n_2306;
assign n_2423 = ~n_2421 & ~n_2422;
assign n_2424 =  x_1975 & ~n_2423;
assign n_2425 = ~x_1975 &  n_2423;
assign n_2426 = ~n_2424 & ~n_2425;
assign n_2427 =  x_1974 & ~n_2306;
assign n_2428 =  i_12 &  n_2306;
assign n_2429 = ~n_2427 & ~n_2428;
assign n_2430 =  x_1974 & ~n_2429;
assign n_2431 = ~x_1974 &  n_2429;
assign n_2432 = ~n_2430 & ~n_2431;
assign n_2433 =  x_1973 & ~n_2306;
assign n_2434 =  i_11 &  n_2306;
assign n_2435 = ~n_2433 & ~n_2434;
assign n_2436 =  x_1973 & ~n_2435;
assign n_2437 = ~x_1973 &  n_2435;
assign n_2438 = ~n_2436 & ~n_2437;
assign n_2439 =  x_1972 & ~n_2306;
assign n_2440 =  i_10 &  n_2306;
assign n_2441 = ~n_2439 & ~n_2440;
assign n_2442 =  x_1972 & ~n_2441;
assign n_2443 = ~x_1972 &  n_2441;
assign n_2444 = ~n_2442 & ~n_2443;
assign n_2445 =  x_1971 & ~n_2306;
assign n_2446 =  i_9 &  n_2306;
assign n_2447 = ~n_2445 & ~n_2446;
assign n_2448 =  x_1971 & ~n_2447;
assign n_2449 = ~x_1971 &  n_2447;
assign n_2450 = ~n_2448 & ~n_2449;
assign n_2451 =  x_1970 & ~n_2306;
assign n_2452 =  i_8 &  n_2306;
assign n_2453 = ~n_2451 & ~n_2452;
assign n_2454 =  x_1970 & ~n_2453;
assign n_2455 = ~x_1970 &  n_2453;
assign n_2456 = ~n_2454 & ~n_2455;
assign n_2457 =  x_1969 & ~n_2306;
assign n_2458 =  i_7 &  n_2306;
assign n_2459 = ~n_2457 & ~n_2458;
assign n_2460 =  x_1969 & ~n_2459;
assign n_2461 = ~x_1969 &  n_2459;
assign n_2462 = ~n_2460 & ~n_2461;
assign n_2463 =  x_1968 & ~n_2306;
assign n_2464 =  i_6 &  n_2306;
assign n_2465 = ~n_2463 & ~n_2464;
assign n_2466 =  x_1968 & ~n_2465;
assign n_2467 = ~x_1968 &  n_2465;
assign n_2468 = ~n_2466 & ~n_2467;
assign n_2469 =  x_1967 & ~n_2306;
assign n_2470 =  i_5 &  n_2306;
assign n_2471 = ~n_2469 & ~n_2470;
assign n_2472 =  x_1967 & ~n_2471;
assign n_2473 = ~x_1967 &  n_2471;
assign n_2474 = ~n_2472 & ~n_2473;
assign n_2475 =  x_1966 & ~n_2306;
assign n_2476 =  i_4 &  n_2306;
assign n_2477 = ~n_2475 & ~n_2476;
assign n_2478 =  x_1966 & ~n_2477;
assign n_2479 = ~x_1966 &  n_2477;
assign n_2480 = ~n_2478 & ~n_2479;
assign n_2481 =  x_1965 & ~n_2306;
assign n_2482 =  i_3 &  n_2306;
assign n_2483 = ~n_2481 & ~n_2482;
assign n_2484 =  x_1965 & ~n_2483;
assign n_2485 = ~x_1965 &  n_2483;
assign n_2486 = ~n_2484 & ~n_2485;
assign n_2487 =  x_1964 & ~n_2306;
assign n_2488 =  i_2 &  n_2306;
assign n_2489 = ~n_2487 & ~n_2488;
assign n_2490 =  x_1964 & ~n_2489;
assign n_2491 = ~x_1964 &  n_2489;
assign n_2492 = ~n_2490 & ~n_2491;
assign n_2493 =  x_1963 & ~n_2306;
assign n_2494 =  i_1 &  n_2306;
assign n_2495 = ~n_2493 & ~n_2494;
assign n_2496 =  x_1963 & ~n_2495;
assign n_2497 = ~x_1963 &  n_2495;
assign n_2498 = ~n_2496 & ~n_2497;
assign n_2499 =  n_1903 &  n_4;
assign n_2500 =  n_186 &  n_2499;
assign n_2501 =  x_1962 & ~n_2500;
assign n_2502 =  i_32 &  n_2500;
assign n_2503 = ~n_2501 & ~n_2502;
assign n_2504 =  x_1962 & ~n_2503;
assign n_2505 = ~x_1962 &  n_2503;
assign n_2506 = ~n_2504 & ~n_2505;
assign n_2507 =  x_1961 & ~n_2500;
assign n_2508 =  i_31 &  n_2500;
assign n_2509 = ~n_2507 & ~n_2508;
assign n_2510 =  x_1961 & ~n_2509;
assign n_2511 = ~x_1961 &  n_2509;
assign n_2512 = ~n_2510 & ~n_2511;
assign n_2513 =  x_1960 & ~n_2500;
assign n_2514 =  i_30 &  n_2500;
assign n_2515 = ~n_2513 & ~n_2514;
assign n_2516 =  x_1960 & ~n_2515;
assign n_2517 = ~x_1960 &  n_2515;
assign n_2518 = ~n_2516 & ~n_2517;
assign n_2519 =  x_1959 & ~n_2500;
assign n_2520 =  i_29 &  n_2500;
assign n_2521 = ~n_2519 & ~n_2520;
assign n_2522 =  x_1959 & ~n_2521;
assign n_2523 = ~x_1959 &  n_2521;
assign n_2524 = ~n_2522 & ~n_2523;
assign n_2525 =  x_1958 & ~n_2500;
assign n_2526 =  i_28 &  n_2500;
assign n_2527 = ~n_2525 & ~n_2526;
assign n_2528 =  x_1958 & ~n_2527;
assign n_2529 = ~x_1958 &  n_2527;
assign n_2530 = ~n_2528 & ~n_2529;
assign n_2531 =  x_1957 & ~n_2500;
assign n_2532 =  i_27 &  n_2500;
assign n_2533 = ~n_2531 & ~n_2532;
assign n_2534 =  x_1957 & ~n_2533;
assign n_2535 = ~x_1957 &  n_2533;
assign n_2536 = ~n_2534 & ~n_2535;
assign n_2537 =  x_1956 & ~n_2500;
assign n_2538 =  i_26 &  n_2500;
assign n_2539 = ~n_2537 & ~n_2538;
assign n_2540 =  x_1956 & ~n_2539;
assign n_2541 = ~x_1956 &  n_2539;
assign n_2542 = ~n_2540 & ~n_2541;
assign n_2543 =  x_1955 & ~n_2500;
assign n_2544 =  i_25 &  n_2500;
assign n_2545 = ~n_2543 & ~n_2544;
assign n_2546 =  x_1955 & ~n_2545;
assign n_2547 = ~x_1955 &  n_2545;
assign n_2548 = ~n_2546 & ~n_2547;
assign n_2549 =  x_1954 & ~n_2500;
assign n_2550 =  i_24 &  n_2500;
assign n_2551 = ~n_2549 & ~n_2550;
assign n_2552 =  x_1954 & ~n_2551;
assign n_2553 = ~x_1954 &  n_2551;
assign n_2554 = ~n_2552 & ~n_2553;
assign n_2555 =  x_1953 & ~n_2500;
assign n_2556 =  i_23 &  n_2500;
assign n_2557 = ~n_2555 & ~n_2556;
assign n_2558 =  x_1953 & ~n_2557;
assign n_2559 = ~x_1953 &  n_2557;
assign n_2560 = ~n_2558 & ~n_2559;
assign n_2561 =  x_1952 & ~n_2500;
assign n_2562 =  i_22 &  n_2500;
assign n_2563 = ~n_2561 & ~n_2562;
assign n_2564 =  x_1952 & ~n_2563;
assign n_2565 = ~x_1952 &  n_2563;
assign n_2566 = ~n_2564 & ~n_2565;
assign n_2567 =  x_1951 & ~n_2500;
assign n_2568 =  i_21 &  n_2500;
assign n_2569 = ~n_2567 & ~n_2568;
assign n_2570 =  x_1951 & ~n_2569;
assign n_2571 = ~x_1951 &  n_2569;
assign n_2572 = ~n_2570 & ~n_2571;
assign n_2573 =  x_1950 & ~n_2500;
assign n_2574 =  i_20 &  n_2500;
assign n_2575 = ~n_2573 & ~n_2574;
assign n_2576 =  x_1950 & ~n_2575;
assign n_2577 = ~x_1950 &  n_2575;
assign n_2578 = ~n_2576 & ~n_2577;
assign n_2579 =  x_1949 & ~n_2500;
assign n_2580 =  i_19 &  n_2500;
assign n_2581 = ~n_2579 & ~n_2580;
assign n_2582 =  x_1949 & ~n_2581;
assign n_2583 = ~x_1949 &  n_2581;
assign n_2584 = ~n_2582 & ~n_2583;
assign n_2585 =  x_1948 & ~n_2500;
assign n_2586 =  i_18 &  n_2500;
assign n_2587 = ~n_2585 & ~n_2586;
assign n_2588 =  x_1948 & ~n_2587;
assign n_2589 = ~x_1948 &  n_2587;
assign n_2590 = ~n_2588 & ~n_2589;
assign n_2591 =  x_1947 & ~n_2500;
assign n_2592 =  i_17 &  n_2500;
assign n_2593 = ~n_2591 & ~n_2592;
assign n_2594 =  x_1947 & ~n_2593;
assign n_2595 = ~x_1947 &  n_2593;
assign n_2596 = ~n_2594 & ~n_2595;
assign n_2597 =  x_1946 & ~n_2500;
assign n_2598 =  i_16 &  n_2500;
assign n_2599 = ~n_2597 & ~n_2598;
assign n_2600 =  x_1946 & ~n_2599;
assign n_2601 = ~x_1946 &  n_2599;
assign n_2602 = ~n_2600 & ~n_2601;
assign n_2603 =  x_1945 & ~n_2500;
assign n_2604 =  i_15 &  n_2500;
assign n_2605 = ~n_2603 & ~n_2604;
assign n_2606 =  x_1945 & ~n_2605;
assign n_2607 = ~x_1945 &  n_2605;
assign n_2608 = ~n_2606 & ~n_2607;
assign n_2609 =  x_1944 & ~n_2500;
assign n_2610 =  i_14 &  n_2500;
assign n_2611 = ~n_2609 & ~n_2610;
assign n_2612 =  x_1944 & ~n_2611;
assign n_2613 = ~x_1944 &  n_2611;
assign n_2614 = ~n_2612 & ~n_2613;
assign n_2615 =  x_1943 & ~n_2500;
assign n_2616 =  i_13 &  n_2500;
assign n_2617 = ~n_2615 & ~n_2616;
assign n_2618 =  x_1943 & ~n_2617;
assign n_2619 = ~x_1943 &  n_2617;
assign n_2620 = ~n_2618 & ~n_2619;
assign n_2621 =  x_1942 & ~n_2500;
assign n_2622 =  i_12 &  n_2500;
assign n_2623 = ~n_2621 & ~n_2622;
assign n_2624 =  x_1942 & ~n_2623;
assign n_2625 = ~x_1942 &  n_2623;
assign n_2626 = ~n_2624 & ~n_2625;
assign n_2627 =  x_1941 & ~n_2500;
assign n_2628 =  i_11 &  n_2500;
assign n_2629 = ~n_2627 & ~n_2628;
assign n_2630 =  x_1941 & ~n_2629;
assign n_2631 = ~x_1941 &  n_2629;
assign n_2632 = ~n_2630 & ~n_2631;
assign n_2633 =  x_1940 & ~n_2500;
assign n_2634 =  i_10 &  n_2500;
assign n_2635 = ~n_2633 & ~n_2634;
assign n_2636 =  x_1940 & ~n_2635;
assign n_2637 = ~x_1940 &  n_2635;
assign n_2638 = ~n_2636 & ~n_2637;
assign n_2639 =  x_1939 & ~n_2500;
assign n_2640 =  i_9 &  n_2500;
assign n_2641 = ~n_2639 & ~n_2640;
assign n_2642 =  x_1939 & ~n_2641;
assign n_2643 = ~x_1939 &  n_2641;
assign n_2644 = ~n_2642 & ~n_2643;
assign n_2645 =  x_1938 & ~n_2500;
assign n_2646 =  i_8 &  n_2500;
assign n_2647 = ~n_2645 & ~n_2646;
assign n_2648 =  x_1938 & ~n_2647;
assign n_2649 = ~x_1938 &  n_2647;
assign n_2650 = ~n_2648 & ~n_2649;
assign n_2651 =  x_1937 & ~n_2500;
assign n_2652 =  i_7 &  n_2500;
assign n_2653 = ~n_2651 & ~n_2652;
assign n_2654 =  x_1937 & ~n_2653;
assign n_2655 = ~x_1937 &  n_2653;
assign n_2656 = ~n_2654 & ~n_2655;
assign n_2657 =  x_1936 & ~n_2500;
assign n_2658 =  i_6 &  n_2500;
assign n_2659 = ~n_2657 & ~n_2658;
assign n_2660 =  x_1936 & ~n_2659;
assign n_2661 = ~x_1936 &  n_2659;
assign n_2662 = ~n_2660 & ~n_2661;
assign n_2663 =  x_1935 & ~n_2500;
assign n_2664 =  i_5 &  n_2500;
assign n_2665 = ~n_2663 & ~n_2664;
assign n_2666 =  x_1935 & ~n_2665;
assign n_2667 = ~x_1935 &  n_2665;
assign n_2668 = ~n_2666 & ~n_2667;
assign n_2669 =  x_1934 & ~n_2500;
assign n_2670 =  i_4 &  n_2500;
assign n_2671 = ~n_2669 & ~n_2670;
assign n_2672 =  x_1934 & ~n_2671;
assign n_2673 = ~x_1934 &  n_2671;
assign n_2674 = ~n_2672 & ~n_2673;
assign n_2675 =  x_1933 & ~n_2500;
assign n_2676 =  i_3 &  n_2500;
assign n_2677 = ~n_2675 & ~n_2676;
assign n_2678 =  x_1933 & ~n_2677;
assign n_2679 = ~x_1933 &  n_2677;
assign n_2680 = ~n_2678 & ~n_2679;
assign n_2681 =  x_1932 & ~n_2500;
assign n_2682 =  i_2 &  n_2500;
assign n_2683 = ~n_2681 & ~n_2682;
assign n_2684 =  x_1932 & ~n_2683;
assign n_2685 = ~x_1932 &  n_2683;
assign n_2686 = ~n_2684 & ~n_2685;
assign n_2687 =  x_1931 & ~n_2500;
assign n_2688 =  i_1 &  n_2500;
assign n_2689 = ~n_2687 & ~n_2688;
assign n_2690 =  x_1931 & ~n_2689;
assign n_2691 = ~x_1931 &  n_2689;
assign n_2692 = ~n_2690 & ~n_2691;
assign n_2693 =  n_8 &  n_186;
assign n_2694 =  x_1930 & ~n_2693;
assign n_2695 =  i_32 &  n_2693;
assign n_2696 = ~n_2694 & ~n_2695;
assign n_2697 =  x_1930 & ~n_2696;
assign n_2698 = ~x_1930 &  n_2696;
assign n_2699 = ~n_2697 & ~n_2698;
assign n_2700 =  x_1929 & ~n_2693;
assign n_2701 =  i_31 &  n_2693;
assign n_2702 = ~n_2700 & ~n_2701;
assign n_2703 =  x_1929 & ~n_2702;
assign n_2704 = ~x_1929 &  n_2702;
assign n_2705 = ~n_2703 & ~n_2704;
assign n_2706 =  x_1928 & ~n_2693;
assign n_2707 =  i_30 &  n_2693;
assign n_2708 = ~n_2706 & ~n_2707;
assign n_2709 =  x_1928 & ~n_2708;
assign n_2710 = ~x_1928 &  n_2708;
assign n_2711 = ~n_2709 & ~n_2710;
assign n_2712 =  x_1927 & ~n_2693;
assign n_2713 =  i_29 &  n_2693;
assign n_2714 = ~n_2712 & ~n_2713;
assign n_2715 =  x_1927 & ~n_2714;
assign n_2716 = ~x_1927 &  n_2714;
assign n_2717 = ~n_2715 & ~n_2716;
assign n_2718 =  x_1926 & ~n_2693;
assign n_2719 =  i_28 &  n_2693;
assign n_2720 = ~n_2718 & ~n_2719;
assign n_2721 =  x_1926 & ~n_2720;
assign n_2722 = ~x_1926 &  n_2720;
assign n_2723 = ~n_2721 & ~n_2722;
assign n_2724 =  x_1925 & ~n_2693;
assign n_2725 =  i_27 &  n_2693;
assign n_2726 = ~n_2724 & ~n_2725;
assign n_2727 =  x_1925 & ~n_2726;
assign n_2728 = ~x_1925 &  n_2726;
assign n_2729 = ~n_2727 & ~n_2728;
assign n_2730 =  x_1924 & ~n_2693;
assign n_2731 =  i_26 &  n_2693;
assign n_2732 = ~n_2730 & ~n_2731;
assign n_2733 =  x_1924 & ~n_2732;
assign n_2734 = ~x_1924 &  n_2732;
assign n_2735 = ~n_2733 & ~n_2734;
assign n_2736 =  x_1923 & ~n_2693;
assign n_2737 =  i_25 &  n_2693;
assign n_2738 = ~n_2736 & ~n_2737;
assign n_2739 =  x_1923 & ~n_2738;
assign n_2740 = ~x_1923 &  n_2738;
assign n_2741 = ~n_2739 & ~n_2740;
assign n_2742 =  x_1922 & ~n_2693;
assign n_2743 =  i_24 &  n_2693;
assign n_2744 = ~n_2742 & ~n_2743;
assign n_2745 =  x_1922 & ~n_2744;
assign n_2746 = ~x_1922 &  n_2744;
assign n_2747 = ~n_2745 & ~n_2746;
assign n_2748 =  x_1921 & ~n_2693;
assign n_2749 =  i_23 &  n_2693;
assign n_2750 = ~n_2748 & ~n_2749;
assign n_2751 =  x_1921 & ~n_2750;
assign n_2752 = ~x_1921 &  n_2750;
assign n_2753 = ~n_2751 & ~n_2752;
assign n_2754 =  x_1920 & ~n_2693;
assign n_2755 =  i_22 &  n_2693;
assign n_2756 = ~n_2754 & ~n_2755;
assign n_2757 =  x_1920 & ~n_2756;
assign n_2758 = ~x_1920 &  n_2756;
assign n_2759 = ~n_2757 & ~n_2758;
assign n_2760 =  x_1919 & ~n_2693;
assign n_2761 =  i_21 &  n_2693;
assign n_2762 = ~n_2760 & ~n_2761;
assign n_2763 =  x_1919 & ~n_2762;
assign n_2764 = ~x_1919 &  n_2762;
assign n_2765 = ~n_2763 & ~n_2764;
assign n_2766 =  x_1918 & ~n_2693;
assign n_2767 =  i_20 &  n_2693;
assign n_2768 = ~n_2766 & ~n_2767;
assign n_2769 =  x_1918 & ~n_2768;
assign n_2770 = ~x_1918 &  n_2768;
assign n_2771 = ~n_2769 & ~n_2770;
assign n_2772 =  x_1917 & ~n_2693;
assign n_2773 =  i_19 &  n_2693;
assign n_2774 = ~n_2772 & ~n_2773;
assign n_2775 =  x_1917 & ~n_2774;
assign n_2776 = ~x_1917 &  n_2774;
assign n_2777 = ~n_2775 & ~n_2776;
assign n_2778 =  x_1916 & ~n_2693;
assign n_2779 =  i_18 &  n_2693;
assign n_2780 = ~n_2778 & ~n_2779;
assign n_2781 =  x_1916 & ~n_2780;
assign n_2782 = ~x_1916 &  n_2780;
assign n_2783 = ~n_2781 & ~n_2782;
assign n_2784 =  x_1915 & ~n_2693;
assign n_2785 =  i_17 &  n_2693;
assign n_2786 = ~n_2784 & ~n_2785;
assign n_2787 =  x_1915 & ~n_2786;
assign n_2788 = ~x_1915 &  n_2786;
assign n_2789 = ~n_2787 & ~n_2788;
assign n_2790 =  x_1914 & ~n_2693;
assign n_2791 =  i_16 &  n_2693;
assign n_2792 = ~n_2790 & ~n_2791;
assign n_2793 =  x_1914 & ~n_2792;
assign n_2794 = ~x_1914 &  n_2792;
assign n_2795 = ~n_2793 & ~n_2794;
assign n_2796 =  x_1913 & ~n_2693;
assign n_2797 =  i_15 &  n_2693;
assign n_2798 = ~n_2796 & ~n_2797;
assign n_2799 =  x_1913 & ~n_2798;
assign n_2800 = ~x_1913 &  n_2798;
assign n_2801 = ~n_2799 & ~n_2800;
assign n_2802 =  x_1912 & ~n_2693;
assign n_2803 =  i_14 &  n_2693;
assign n_2804 = ~n_2802 & ~n_2803;
assign n_2805 =  x_1912 & ~n_2804;
assign n_2806 = ~x_1912 &  n_2804;
assign n_2807 = ~n_2805 & ~n_2806;
assign n_2808 =  x_1911 & ~n_2693;
assign n_2809 =  i_13 &  n_2693;
assign n_2810 = ~n_2808 & ~n_2809;
assign n_2811 =  x_1911 & ~n_2810;
assign n_2812 = ~x_1911 &  n_2810;
assign n_2813 = ~n_2811 & ~n_2812;
assign n_2814 =  x_1910 & ~n_2693;
assign n_2815 =  i_12 &  n_2693;
assign n_2816 = ~n_2814 & ~n_2815;
assign n_2817 =  x_1910 & ~n_2816;
assign n_2818 = ~x_1910 &  n_2816;
assign n_2819 = ~n_2817 & ~n_2818;
assign n_2820 =  x_1909 & ~n_2693;
assign n_2821 =  i_11 &  n_2693;
assign n_2822 = ~n_2820 & ~n_2821;
assign n_2823 =  x_1909 & ~n_2822;
assign n_2824 = ~x_1909 &  n_2822;
assign n_2825 = ~n_2823 & ~n_2824;
assign n_2826 =  x_1908 & ~n_2693;
assign n_2827 =  i_10 &  n_2693;
assign n_2828 = ~n_2826 & ~n_2827;
assign n_2829 =  x_1908 & ~n_2828;
assign n_2830 = ~x_1908 &  n_2828;
assign n_2831 = ~n_2829 & ~n_2830;
assign n_2832 =  x_1907 & ~n_2693;
assign n_2833 =  i_9 &  n_2693;
assign n_2834 = ~n_2832 & ~n_2833;
assign n_2835 =  x_1907 & ~n_2834;
assign n_2836 = ~x_1907 &  n_2834;
assign n_2837 = ~n_2835 & ~n_2836;
assign n_2838 =  x_1906 & ~n_2693;
assign n_2839 =  i_8 &  n_2693;
assign n_2840 = ~n_2838 & ~n_2839;
assign n_2841 =  x_1906 & ~n_2840;
assign n_2842 = ~x_1906 &  n_2840;
assign n_2843 = ~n_2841 & ~n_2842;
assign n_2844 =  x_1905 & ~n_2693;
assign n_2845 =  i_7 &  n_2693;
assign n_2846 = ~n_2844 & ~n_2845;
assign n_2847 =  x_1905 & ~n_2846;
assign n_2848 = ~x_1905 &  n_2846;
assign n_2849 = ~n_2847 & ~n_2848;
assign n_2850 =  x_1904 & ~n_2693;
assign n_2851 =  i_6 &  n_2693;
assign n_2852 = ~n_2850 & ~n_2851;
assign n_2853 =  x_1904 & ~n_2852;
assign n_2854 = ~x_1904 &  n_2852;
assign n_2855 = ~n_2853 & ~n_2854;
assign n_2856 =  x_1903 & ~n_2693;
assign n_2857 =  i_5 &  n_2693;
assign n_2858 = ~n_2856 & ~n_2857;
assign n_2859 =  x_1903 & ~n_2858;
assign n_2860 = ~x_1903 &  n_2858;
assign n_2861 = ~n_2859 & ~n_2860;
assign n_2862 =  x_1902 & ~n_2693;
assign n_2863 =  i_4 &  n_2693;
assign n_2864 = ~n_2862 & ~n_2863;
assign n_2865 =  x_1902 & ~n_2864;
assign n_2866 = ~x_1902 &  n_2864;
assign n_2867 = ~n_2865 & ~n_2866;
assign n_2868 =  x_1901 & ~n_2693;
assign n_2869 =  i_3 &  n_2693;
assign n_2870 = ~n_2868 & ~n_2869;
assign n_2871 =  x_1901 & ~n_2870;
assign n_2872 = ~x_1901 &  n_2870;
assign n_2873 = ~n_2871 & ~n_2872;
assign n_2874 =  x_1900 & ~n_2693;
assign n_2875 =  i_2 &  n_2693;
assign n_2876 = ~n_2874 & ~n_2875;
assign n_2877 =  x_1900 & ~n_2876;
assign n_2878 = ~x_1900 &  n_2876;
assign n_2879 = ~n_2877 & ~n_2878;
assign n_2880 =  x_1899 & ~n_2693;
assign n_2881 =  i_1 &  n_2693;
assign n_2882 = ~n_2880 & ~n_2881;
assign n_2883 =  x_1899 & ~n_2882;
assign n_2884 = ~x_1899 &  n_2882;
assign n_2885 = ~n_2883 & ~n_2884;
assign n_2886 =  x_38 & ~x_39;
assign n_2887 =  n_586 &  n_2886;
assign n_2888 =  n_2296 &  n_2887;
assign n_2889 =  x_1898 & ~n_2888;
assign n_2890 =  i_32 &  n_2888;
assign n_2891 = ~n_2889 & ~n_2890;
assign n_2892 =  x_1898 & ~n_2891;
assign n_2893 = ~x_1898 &  n_2891;
assign n_2894 = ~n_2892 & ~n_2893;
assign n_2895 =  x_1897 & ~n_2888;
assign n_2896 =  i_31 &  n_2888;
assign n_2897 = ~n_2895 & ~n_2896;
assign n_2898 =  x_1897 & ~n_2897;
assign n_2899 = ~x_1897 &  n_2897;
assign n_2900 = ~n_2898 & ~n_2899;
assign n_2901 =  x_1896 & ~n_2888;
assign n_2902 =  i_30 &  n_2888;
assign n_2903 = ~n_2901 & ~n_2902;
assign n_2904 =  x_1896 & ~n_2903;
assign n_2905 = ~x_1896 &  n_2903;
assign n_2906 = ~n_2904 & ~n_2905;
assign n_2907 =  x_1895 & ~n_2888;
assign n_2908 =  i_29 &  n_2888;
assign n_2909 = ~n_2907 & ~n_2908;
assign n_2910 =  x_1895 & ~n_2909;
assign n_2911 = ~x_1895 &  n_2909;
assign n_2912 = ~n_2910 & ~n_2911;
assign n_2913 =  x_1894 & ~n_2888;
assign n_2914 =  i_28 &  n_2888;
assign n_2915 = ~n_2913 & ~n_2914;
assign n_2916 =  x_1894 & ~n_2915;
assign n_2917 = ~x_1894 &  n_2915;
assign n_2918 = ~n_2916 & ~n_2917;
assign n_2919 =  x_1893 & ~n_2888;
assign n_2920 =  i_27 &  n_2888;
assign n_2921 = ~n_2919 & ~n_2920;
assign n_2922 =  x_1893 & ~n_2921;
assign n_2923 = ~x_1893 &  n_2921;
assign n_2924 = ~n_2922 & ~n_2923;
assign n_2925 =  x_1892 & ~n_2888;
assign n_2926 =  i_26 &  n_2888;
assign n_2927 = ~n_2925 & ~n_2926;
assign n_2928 =  x_1892 & ~n_2927;
assign n_2929 = ~x_1892 &  n_2927;
assign n_2930 = ~n_2928 & ~n_2929;
assign n_2931 =  x_1891 & ~n_2888;
assign n_2932 =  i_25 &  n_2888;
assign n_2933 = ~n_2931 & ~n_2932;
assign n_2934 =  x_1891 & ~n_2933;
assign n_2935 = ~x_1891 &  n_2933;
assign n_2936 = ~n_2934 & ~n_2935;
assign n_2937 =  x_1890 & ~n_2888;
assign n_2938 =  i_24 &  n_2888;
assign n_2939 = ~n_2937 & ~n_2938;
assign n_2940 =  x_1890 & ~n_2939;
assign n_2941 = ~x_1890 &  n_2939;
assign n_2942 = ~n_2940 & ~n_2941;
assign n_2943 =  x_1889 & ~n_2888;
assign n_2944 =  i_23 &  n_2888;
assign n_2945 = ~n_2943 & ~n_2944;
assign n_2946 =  x_1889 & ~n_2945;
assign n_2947 = ~x_1889 &  n_2945;
assign n_2948 = ~n_2946 & ~n_2947;
assign n_2949 =  x_1888 & ~n_2888;
assign n_2950 =  i_22 &  n_2888;
assign n_2951 = ~n_2949 & ~n_2950;
assign n_2952 =  x_1888 & ~n_2951;
assign n_2953 = ~x_1888 &  n_2951;
assign n_2954 = ~n_2952 & ~n_2953;
assign n_2955 =  x_1887 & ~n_2888;
assign n_2956 =  i_21 &  n_2888;
assign n_2957 = ~n_2955 & ~n_2956;
assign n_2958 =  x_1887 & ~n_2957;
assign n_2959 = ~x_1887 &  n_2957;
assign n_2960 = ~n_2958 & ~n_2959;
assign n_2961 =  x_1886 & ~n_2888;
assign n_2962 =  i_20 &  n_2888;
assign n_2963 = ~n_2961 & ~n_2962;
assign n_2964 =  x_1886 & ~n_2963;
assign n_2965 = ~x_1886 &  n_2963;
assign n_2966 = ~n_2964 & ~n_2965;
assign n_2967 =  x_1885 & ~n_2888;
assign n_2968 =  i_19 &  n_2888;
assign n_2969 = ~n_2967 & ~n_2968;
assign n_2970 =  x_1885 & ~n_2969;
assign n_2971 = ~x_1885 &  n_2969;
assign n_2972 = ~n_2970 & ~n_2971;
assign n_2973 =  x_1884 & ~n_2888;
assign n_2974 =  i_18 &  n_2888;
assign n_2975 = ~n_2973 & ~n_2974;
assign n_2976 =  x_1884 & ~n_2975;
assign n_2977 = ~x_1884 &  n_2975;
assign n_2978 = ~n_2976 & ~n_2977;
assign n_2979 =  x_1883 & ~n_2888;
assign n_2980 =  i_17 &  n_2888;
assign n_2981 = ~n_2979 & ~n_2980;
assign n_2982 =  x_1883 & ~n_2981;
assign n_2983 = ~x_1883 &  n_2981;
assign n_2984 = ~n_2982 & ~n_2983;
assign n_2985 =  x_1882 & ~n_2888;
assign n_2986 =  i_16 &  n_2888;
assign n_2987 = ~n_2985 & ~n_2986;
assign n_2988 =  x_1882 & ~n_2987;
assign n_2989 = ~x_1882 &  n_2987;
assign n_2990 = ~n_2988 & ~n_2989;
assign n_2991 =  x_1881 & ~n_2888;
assign n_2992 =  i_15 &  n_2888;
assign n_2993 = ~n_2991 & ~n_2992;
assign n_2994 =  x_1881 & ~n_2993;
assign n_2995 = ~x_1881 &  n_2993;
assign n_2996 = ~n_2994 & ~n_2995;
assign n_2997 =  x_1880 & ~n_2888;
assign n_2998 =  i_14 &  n_2888;
assign n_2999 = ~n_2997 & ~n_2998;
assign n_3000 =  x_1880 & ~n_2999;
assign n_3001 = ~x_1880 &  n_2999;
assign n_3002 = ~n_3000 & ~n_3001;
assign n_3003 =  x_1879 & ~n_2888;
assign n_3004 =  i_13 &  n_2888;
assign n_3005 = ~n_3003 & ~n_3004;
assign n_3006 =  x_1879 & ~n_3005;
assign n_3007 = ~x_1879 &  n_3005;
assign n_3008 = ~n_3006 & ~n_3007;
assign n_3009 =  x_1878 & ~n_2888;
assign n_3010 =  i_12 &  n_2888;
assign n_3011 = ~n_3009 & ~n_3010;
assign n_3012 =  x_1878 & ~n_3011;
assign n_3013 = ~x_1878 &  n_3011;
assign n_3014 = ~n_3012 & ~n_3013;
assign n_3015 =  x_1877 & ~n_2888;
assign n_3016 =  i_11 &  n_2888;
assign n_3017 = ~n_3015 & ~n_3016;
assign n_3018 =  x_1877 & ~n_3017;
assign n_3019 = ~x_1877 &  n_3017;
assign n_3020 = ~n_3018 & ~n_3019;
assign n_3021 =  x_1876 & ~n_2888;
assign n_3022 =  i_10 &  n_2888;
assign n_3023 = ~n_3021 & ~n_3022;
assign n_3024 =  x_1876 & ~n_3023;
assign n_3025 = ~x_1876 &  n_3023;
assign n_3026 = ~n_3024 & ~n_3025;
assign n_3027 =  x_1875 & ~n_2888;
assign n_3028 =  i_9 &  n_2888;
assign n_3029 = ~n_3027 & ~n_3028;
assign n_3030 =  x_1875 & ~n_3029;
assign n_3031 = ~x_1875 &  n_3029;
assign n_3032 = ~n_3030 & ~n_3031;
assign n_3033 =  x_1874 & ~n_2888;
assign n_3034 =  i_8 &  n_2888;
assign n_3035 = ~n_3033 & ~n_3034;
assign n_3036 =  x_1874 & ~n_3035;
assign n_3037 = ~x_1874 &  n_3035;
assign n_3038 = ~n_3036 & ~n_3037;
assign n_3039 =  x_1873 & ~n_2888;
assign n_3040 =  i_7 &  n_2888;
assign n_3041 = ~n_3039 & ~n_3040;
assign n_3042 =  x_1873 & ~n_3041;
assign n_3043 = ~x_1873 &  n_3041;
assign n_3044 = ~n_3042 & ~n_3043;
assign n_3045 =  x_1872 & ~n_2888;
assign n_3046 =  i_6 &  n_2888;
assign n_3047 = ~n_3045 & ~n_3046;
assign n_3048 =  x_1872 & ~n_3047;
assign n_3049 = ~x_1872 &  n_3047;
assign n_3050 = ~n_3048 & ~n_3049;
assign n_3051 =  x_1871 & ~n_2888;
assign n_3052 =  i_5 &  n_2888;
assign n_3053 = ~n_3051 & ~n_3052;
assign n_3054 =  x_1871 & ~n_3053;
assign n_3055 = ~x_1871 &  n_3053;
assign n_3056 = ~n_3054 & ~n_3055;
assign n_3057 =  x_1870 & ~n_2888;
assign n_3058 =  i_4 &  n_2888;
assign n_3059 = ~n_3057 & ~n_3058;
assign n_3060 =  x_1870 & ~n_3059;
assign n_3061 = ~x_1870 &  n_3059;
assign n_3062 = ~n_3060 & ~n_3061;
assign n_3063 =  x_1869 & ~n_2888;
assign n_3064 =  i_3 &  n_2888;
assign n_3065 = ~n_3063 & ~n_3064;
assign n_3066 =  x_1869 & ~n_3065;
assign n_3067 = ~x_1869 &  n_3065;
assign n_3068 = ~n_3066 & ~n_3067;
assign n_3069 =  x_1868 & ~n_2888;
assign n_3070 =  i_2 &  n_2888;
assign n_3071 = ~n_3069 & ~n_3070;
assign n_3072 =  x_1868 & ~n_3071;
assign n_3073 = ~x_1868 &  n_3071;
assign n_3074 = ~n_3072 & ~n_3073;
assign n_3075 =  x_1867 & ~n_2888;
assign n_3076 =  i_1 &  n_2888;
assign n_3077 = ~n_3075 & ~n_3076;
assign n_3078 =  x_1867 & ~n_3077;
assign n_3079 = ~x_1867 &  n_3077;
assign n_3080 = ~n_3078 & ~n_3079;
assign n_3081 =  n_1708 &  n_4;
assign n_3082 =  n_3081 &  n_186;
assign n_3083 =  x_1866 & ~n_3082;
assign n_3084 =  i_32 &  n_3082;
assign n_3085 = ~n_3083 & ~n_3084;
assign n_3086 =  x_1866 & ~n_3085;
assign n_3087 = ~x_1866 &  n_3085;
assign n_3088 = ~n_3086 & ~n_3087;
assign n_3089 =  x_1865 & ~n_3082;
assign n_3090 =  i_31 &  n_3082;
assign n_3091 = ~n_3089 & ~n_3090;
assign n_3092 =  x_1865 & ~n_3091;
assign n_3093 = ~x_1865 &  n_3091;
assign n_3094 = ~n_3092 & ~n_3093;
assign n_3095 =  x_1864 & ~n_3082;
assign n_3096 =  i_30 &  n_3082;
assign n_3097 = ~n_3095 & ~n_3096;
assign n_3098 =  x_1864 & ~n_3097;
assign n_3099 = ~x_1864 &  n_3097;
assign n_3100 = ~n_3098 & ~n_3099;
assign n_3101 =  x_1863 & ~n_3082;
assign n_3102 =  i_29 &  n_3082;
assign n_3103 = ~n_3101 & ~n_3102;
assign n_3104 =  x_1863 & ~n_3103;
assign n_3105 = ~x_1863 &  n_3103;
assign n_3106 = ~n_3104 & ~n_3105;
assign n_3107 =  x_1862 & ~n_3082;
assign n_3108 =  i_28 &  n_3082;
assign n_3109 = ~n_3107 & ~n_3108;
assign n_3110 =  x_1862 & ~n_3109;
assign n_3111 = ~x_1862 &  n_3109;
assign n_3112 = ~n_3110 & ~n_3111;
assign n_3113 =  x_1861 & ~n_3082;
assign n_3114 =  i_27 &  n_3082;
assign n_3115 = ~n_3113 & ~n_3114;
assign n_3116 =  x_1861 & ~n_3115;
assign n_3117 = ~x_1861 &  n_3115;
assign n_3118 = ~n_3116 & ~n_3117;
assign n_3119 =  x_1860 & ~n_3082;
assign n_3120 =  i_26 &  n_3082;
assign n_3121 = ~n_3119 & ~n_3120;
assign n_3122 =  x_1860 & ~n_3121;
assign n_3123 = ~x_1860 &  n_3121;
assign n_3124 = ~n_3122 & ~n_3123;
assign n_3125 =  x_1859 & ~n_3082;
assign n_3126 =  i_25 &  n_3082;
assign n_3127 = ~n_3125 & ~n_3126;
assign n_3128 =  x_1859 & ~n_3127;
assign n_3129 = ~x_1859 &  n_3127;
assign n_3130 = ~n_3128 & ~n_3129;
assign n_3131 =  x_1858 & ~n_3082;
assign n_3132 =  i_24 &  n_3082;
assign n_3133 = ~n_3131 & ~n_3132;
assign n_3134 =  x_1858 & ~n_3133;
assign n_3135 = ~x_1858 &  n_3133;
assign n_3136 = ~n_3134 & ~n_3135;
assign n_3137 =  x_1857 & ~n_3082;
assign n_3138 =  i_23 &  n_3082;
assign n_3139 = ~n_3137 & ~n_3138;
assign n_3140 =  x_1857 & ~n_3139;
assign n_3141 = ~x_1857 &  n_3139;
assign n_3142 = ~n_3140 & ~n_3141;
assign n_3143 =  x_1856 & ~n_3082;
assign n_3144 =  i_22 &  n_3082;
assign n_3145 = ~n_3143 & ~n_3144;
assign n_3146 =  x_1856 & ~n_3145;
assign n_3147 = ~x_1856 &  n_3145;
assign n_3148 = ~n_3146 & ~n_3147;
assign n_3149 =  x_1855 & ~n_3082;
assign n_3150 =  i_21 &  n_3082;
assign n_3151 = ~n_3149 & ~n_3150;
assign n_3152 =  x_1855 & ~n_3151;
assign n_3153 = ~x_1855 &  n_3151;
assign n_3154 = ~n_3152 & ~n_3153;
assign n_3155 =  x_1854 & ~n_3082;
assign n_3156 =  i_20 &  n_3082;
assign n_3157 = ~n_3155 & ~n_3156;
assign n_3158 =  x_1854 & ~n_3157;
assign n_3159 = ~x_1854 &  n_3157;
assign n_3160 = ~n_3158 & ~n_3159;
assign n_3161 =  x_1853 & ~n_3082;
assign n_3162 =  i_19 &  n_3082;
assign n_3163 = ~n_3161 & ~n_3162;
assign n_3164 =  x_1853 & ~n_3163;
assign n_3165 = ~x_1853 &  n_3163;
assign n_3166 = ~n_3164 & ~n_3165;
assign n_3167 =  x_1852 & ~n_3082;
assign n_3168 =  i_18 &  n_3082;
assign n_3169 = ~n_3167 & ~n_3168;
assign n_3170 =  x_1852 & ~n_3169;
assign n_3171 = ~x_1852 &  n_3169;
assign n_3172 = ~n_3170 & ~n_3171;
assign n_3173 =  x_1851 & ~n_3082;
assign n_3174 =  i_17 &  n_3082;
assign n_3175 = ~n_3173 & ~n_3174;
assign n_3176 =  x_1851 & ~n_3175;
assign n_3177 = ~x_1851 &  n_3175;
assign n_3178 = ~n_3176 & ~n_3177;
assign n_3179 =  x_1850 & ~n_3082;
assign n_3180 =  i_16 &  n_3082;
assign n_3181 = ~n_3179 & ~n_3180;
assign n_3182 =  x_1850 & ~n_3181;
assign n_3183 = ~x_1850 &  n_3181;
assign n_3184 = ~n_3182 & ~n_3183;
assign n_3185 =  x_1849 & ~n_3082;
assign n_3186 =  i_15 &  n_3082;
assign n_3187 = ~n_3185 & ~n_3186;
assign n_3188 =  x_1849 & ~n_3187;
assign n_3189 = ~x_1849 &  n_3187;
assign n_3190 = ~n_3188 & ~n_3189;
assign n_3191 =  x_1848 & ~n_3082;
assign n_3192 =  i_14 &  n_3082;
assign n_3193 = ~n_3191 & ~n_3192;
assign n_3194 =  x_1848 & ~n_3193;
assign n_3195 = ~x_1848 &  n_3193;
assign n_3196 = ~n_3194 & ~n_3195;
assign n_3197 =  x_1847 & ~n_3082;
assign n_3198 =  i_13 &  n_3082;
assign n_3199 = ~n_3197 & ~n_3198;
assign n_3200 =  x_1847 & ~n_3199;
assign n_3201 = ~x_1847 &  n_3199;
assign n_3202 = ~n_3200 & ~n_3201;
assign n_3203 =  x_1846 & ~n_3082;
assign n_3204 =  i_12 &  n_3082;
assign n_3205 = ~n_3203 & ~n_3204;
assign n_3206 =  x_1846 & ~n_3205;
assign n_3207 = ~x_1846 &  n_3205;
assign n_3208 = ~n_3206 & ~n_3207;
assign n_3209 =  x_1845 & ~n_3082;
assign n_3210 =  i_11 &  n_3082;
assign n_3211 = ~n_3209 & ~n_3210;
assign n_3212 =  x_1845 & ~n_3211;
assign n_3213 = ~x_1845 &  n_3211;
assign n_3214 = ~n_3212 & ~n_3213;
assign n_3215 =  x_1844 & ~n_3082;
assign n_3216 =  i_10 &  n_3082;
assign n_3217 = ~n_3215 & ~n_3216;
assign n_3218 =  x_1844 & ~n_3217;
assign n_3219 = ~x_1844 &  n_3217;
assign n_3220 = ~n_3218 & ~n_3219;
assign n_3221 =  x_1843 & ~n_3082;
assign n_3222 =  i_9 &  n_3082;
assign n_3223 = ~n_3221 & ~n_3222;
assign n_3224 =  x_1843 & ~n_3223;
assign n_3225 = ~x_1843 &  n_3223;
assign n_3226 = ~n_3224 & ~n_3225;
assign n_3227 =  x_1842 & ~n_3082;
assign n_3228 =  i_8 &  n_3082;
assign n_3229 = ~n_3227 & ~n_3228;
assign n_3230 =  x_1842 & ~n_3229;
assign n_3231 = ~x_1842 &  n_3229;
assign n_3232 = ~n_3230 & ~n_3231;
assign n_3233 =  x_1841 & ~n_3082;
assign n_3234 =  i_7 &  n_3082;
assign n_3235 = ~n_3233 & ~n_3234;
assign n_3236 =  x_1841 & ~n_3235;
assign n_3237 = ~x_1841 &  n_3235;
assign n_3238 = ~n_3236 & ~n_3237;
assign n_3239 =  x_1840 & ~n_3082;
assign n_3240 =  i_6 &  n_3082;
assign n_3241 = ~n_3239 & ~n_3240;
assign n_3242 =  x_1840 & ~n_3241;
assign n_3243 = ~x_1840 &  n_3241;
assign n_3244 = ~n_3242 & ~n_3243;
assign n_3245 =  x_1839 & ~n_3082;
assign n_3246 =  i_5 &  n_3082;
assign n_3247 = ~n_3245 & ~n_3246;
assign n_3248 =  x_1839 & ~n_3247;
assign n_3249 = ~x_1839 &  n_3247;
assign n_3250 = ~n_3248 & ~n_3249;
assign n_3251 =  x_1838 & ~n_3082;
assign n_3252 =  i_4 &  n_3082;
assign n_3253 = ~n_3251 & ~n_3252;
assign n_3254 =  x_1838 & ~n_3253;
assign n_3255 = ~x_1838 &  n_3253;
assign n_3256 = ~n_3254 & ~n_3255;
assign n_3257 =  x_1837 & ~n_3082;
assign n_3258 =  i_3 &  n_3082;
assign n_3259 = ~n_3257 & ~n_3258;
assign n_3260 =  x_1837 & ~n_3259;
assign n_3261 = ~x_1837 &  n_3259;
assign n_3262 = ~n_3260 & ~n_3261;
assign n_3263 =  x_1836 & ~n_3082;
assign n_3264 =  i_2 &  n_3082;
assign n_3265 = ~n_3263 & ~n_3264;
assign n_3266 =  x_1836 & ~n_3265;
assign n_3267 = ~x_1836 &  n_3265;
assign n_3268 = ~n_3266 & ~n_3267;
assign n_3269 =  x_1835 & ~n_3082;
assign n_3270 =  i_1 &  n_3082;
assign n_3271 = ~n_3269 & ~n_3270;
assign n_3272 =  x_1835 & ~n_3271;
assign n_3273 = ~x_1835 &  n_3271;
assign n_3274 = ~n_3272 & ~n_3273;
assign n_3275 =  n_190 &  n_4;
assign n_3276 =  n_186 &  n_3275;
assign n_3277 =  x_1834 & ~n_3276;
assign n_3278 =  i_32 &  n_3276;
assign n_3279 = ~n_3277 & ~n_3278;
assign n_3280 =  x_1834 & ~n_3279;
assign n_3281 = ~x_1834 &  n_3279;
assign n_3282 = ~n_3280 & ~n_3281;
assign n_3283 =  x_1833 & ~n_3276;
assign n_3284 =  i_31 &  n_3276;
assign n_3285 = ~n_3283 & ~n_3284;
assign n_3286 =  x_1833 & ~n_3285;
assign n_3287 = ~x_1833 &  n_3285;
assign n_3288 = ~n_3286 & ~n_3287;
assign n_3289 =  x_1832 & ~n_3276;
assign n_3290 =  i_30 &  n_3276;
assign n_3291 = ~n_3289 & ~n_3290;
assign n_3292 =  x_1832 & ~n_3291;
assign n_3293 = ~x_1832 &  n_3291;
assign n_3294 = ~n_3292 & ~n_3293;
assign n_3295 =  x_1831 & ~n_3276;
assign n_3296 =  i_29 &  n_3276;
assign n_3297 = ~n_3295 & ~n_3296;
assign n_3298 =  x_1831 & ~n_3297;
assign n_3299 = ~x_1831 &  n_3297;
assign n_3300 = ~n_3298 & ~n_3299;
assign n_3301 =  x_1830 & ~n_3276;
assign n_3302 =  i_28 &  n_3276;
assign n_3303 = ~n_3301 & ~n_3302;
assign n_3304 =  x_1830 & ~n_3303;
assign n_3305 = ~x_1830 &  n_3303;
assign n_3306 = ~n_3304 & ~n_3305;
assign n_3307 =  x_1829 & ~n_3276;
assign n_3308 =  i_27 &  n_3276;
assign n_3309 = ~n_3307 & ~n_3308;
assign n_3310 =  x_1829 & ~n_3309;
assign n_3311 = ~x_1829 &  n_3309;
assign n_3312 = ~n_3310 & ~n_3311;
assign n_3313 =  x_1828 & ~n_3276;
assign n_3314 =  i_26 &  n_3276;
assign n_3315 = ~n_3313 & ~n_3314;
assign n_3316 =  x_1828 & ~n_3315;
assign n_3317 = ~x_1828 &  n_3315;
assign n_3318 = ~n_3316 & ~n_3317;
assign n_3319 =  x_1827 & ~n_3276;
assign n_3320 =  i_25 &  n_3276;
assign n_3321 = ~n_3319 & ~n_3320;
assign n_3322 =  x_1827 & ~n_3321;
assign n_3323 = ~x_1827 &  n_3321;
assign n_3324 = ~n_3322 & ~n_3323;
assign n_3325 =  x_1826 & ~n_3276;
assign n_3326 =  i_24 &  n_3276;
assign n_3327 = ~n_3325 & ~n_3326;
assign n_3328 =  x_1826 & ~n_3327;
assign n_3329 = ~x_1826 &  n_3327;
assign n_3330 = ~n_3328 & ~n_3329;
assign n_3331 =  x_1825 & ~n_3276;
assign n_3332 =  i_23 &  n_3276;
assign n_3333 = ~n_3331 & ~n_3332;
assign n_3334 =  x_1825 & ~n_3333;
assign n_3335 = ~x_1825 &  n_3333;
assign n_3336 = ~n_3334 & ~n_3335;
assign n_3337 =  x_1824 & ~n_3276;
assign n_3338 =  i_22 &  n_3276;
assign n_3339 = ~n_3337 & ~n_3338;
assign n_3340 =  x_1824 & ~n_3339;
assign n_3341 = ~x_1824 &  n_3339;
assign n_3342 = ~n_3340 & ~n_3341;
assign n_3343 =  x_1823 & ~n_3276;
assign n_3344 =  i_21 &  n_3276;
assign n_3345 = ~n_3343 & ~n_3344;
assign n_3346 =  x_1823 & ~n_3345;
assign n_3347 = ~x_1823 &  n_3345;
assign n_3348 = ~n_3346 & ~n_3347;
assign n_3349 =  x_1822 & ~n_3276;
assign n_3350 =  i_20 &  n_3276;
assign n_3351 = ~n_3349 & ~n_3350;
assign n_3352 =  x_1822 & ~n_3351;
assign n_3353 = ~x_1822 &  n_3351;
assign n_3354 = ~n_3352 & ~n_3353;
assign n_3355 =  x_1821 & ~n_3276;
assign n_3356 =  i_19 &  n_3276;
assign n_3357 = ~n_3355 & ~n_3356;
assign n_3358 =  x_1821 & ~n_3357;
assign n_3359 = ~x_1821 &  n_3357;
assign n_3360 = ~n_3358 & ~n_3359;
assign n_3361 =  x_1820 & ~n_3276;
assign n_3362 =  i_18 &  n_3276;
assign n_3363 = ~n_3361 & ~n_3362;
assign n_3364 =  x_1820 & ~n_3363;
assign n_3365 = ~x_1820 &  n_3363;
assign n_3366 = ~n_3364 & ~n_3365;
assign n_3367 =  x_1819 & ~n_3276;
assign n_3368 =  i_17 &  n_3276;
assign n_3369 = ~n_3367 & ~n_3368;
assign n_3370 =  x_1819 & ~n_3369;
assign n_3371 = ~x_1819 &  n_3369;
assign n_3372 = ~n_3370 & ~n_3371;
assign n_3373 =  x_1818 & ~n_3276;
assign n_3374 =  i_16 &  n_3276;
assign n_3375 = ~n_3373 & ~n_3374;
assign n_3376 =  x_1818 & ~n_3375;
assign n_3377 = ~x_1818 &  n_3375;
assign n_3378 = ~n_3376 & ~n_3377;
assign n_3379 =  x_1817 & ~n_3276;
assign n_3380 =  i_15 &  n_3276;
assign n_3381 = ~n_3379 & ~n_3380;
assign n_3382 =  x_1817 & ~n_3381;
assign n_3383 = ~x_1817 &  n_3381;
assign n_3384 = ~n_3382 & ~n_3383;
assign n_3385 =  x_1816 & ~n_3276;
assign n_3386 =  i_14 &  n_3276;
assign n_3387 = ~n_3385 & ~n_3386;
assign n_3388 =  x_1816 & ~n_3387;
assign n_3389 = ~x_1816 &  n_3387;
assign n_3390 = ~n_3388 & ~n_3389;
assign n_3391 =  x_1815 & ~n_3276;
assign n_3392 =  i_13 &  n_3276;
assign n_3393 = ~n_3391 & ~n_3392;
assign n_3394 =  x_1815 & ~n_3393;
assign n_3395 = ~x_1815 &  n_3393;
assign n_3396 = ~n_3394 & ~n_3395;
assign n_3397 =  x_1814 & ~n_3276;
assign n_3398 =  i_12 &  n_3276;
assign n_3399 = ~n_3397 & ~n_3398;
assign n_3400 =  x_1814 & ~n_3399;
assign n_3401 = ~x_1814 &  n_3399;
assign n_3402 = ~n_3400 & ~n_3401;
assign n_3403 =  x_1813 & ~n_3276;
assign n_3404 =  i_11 &  n_3276;
assign n_3405 = ~n_3403 & ~n_3404;
assign n_3406 =  x_1813 & ~n_3405;
assign n_3407 = ~x_1813 &  n_3405;
assign n_3408 = ~n_3406 & ~n_3407;
assign n_3409 =  x_1812 & ~n_3276;
assign n_3410 =  i_10 &  n_3276;
assign n_3411 = ~n_3409 & ~n_3410;
assign n_3412 =  x_1812 & ~n_3411;
assign n_3413 = ~x_1812 &  n_3411;
assign n_3414 = ~n_3412 & ~n_3413;
assign n_3415 =  x_1811 & ~n_3276;
assign n_3416 =  i_9 &  n_3276;
assign n_3417 = ~n_3415 & ~n_3416;
assign n_3418 =  x_1811 & ~n_3417;
assign n_3419 = ~x_1811 &  n_3417;
assign n_3420 = ~n_3418 & ~n_3419;
assign n_3421 =  x_1810 & ~n_3276;
assign n_3422 =  i_8 &  n_3276;
assign n_3423 = ~n_3421 & ~n_3422;
assign n_3424 =  x_1810 & ~n_3423;
assign n_3425 = ~x_1810 &  n_3423;
assign n_3426 = ~n_3424 & ~n_3425;
assign n_3427 =  x_1809 & ~n_3276;
assign n_3428 =  i_7 &  n_3276;
assign n_3429 = ~n_3427 & ~n_3428;
assign n_3430 =  x_1809 & ~n_3429;
assign n_3431 = ~x_1809 &  n_3429;
assign n_3432 = ~n_3430 & ~n_3431;
assign n_3433 =  x_1808 & ~n_3276;
assign n_3434 =  i_6 &  n_3276;
assign n_3435 = ~n_3433 & ~n_3434;
assign n_3436 =  x_1808 & ~n_3435;
assign n_3437 = ~x_1808 &  n_3435;
assign n_3438 = ~n_3436 & ~n_3437;
assign n_3439 =  x_1807 & ~n_3276;
assign n_3440 =  i_5 &  n_3276;
assign n_3441 = ~n_3439 & ~n_3440;
assign n_3442 =  x_1807 & ~n_3441;
assign n_3443 = ~x_1807 &  n_3441;
assign n_3444 = ~n_3442 & ~n_3443;
assign n_3445 =  x_1806 & ~n_3276;
assign n_3446 =  i_4 &  n_3276;
assign n_3447 = ~n_3445 & ~n_3446;
assign n_3448 =  x_1806 & ~n_3447;
assign n_3449 = ~x_1806 &  n_3447;
assign n_3450 = ~n_3448 & ~n_3449;
assign n_3451 =  x_1805 & ~n_3276;
assign n_3452 =  i_3 &  n_3276;
assign n_3453 = ~n_3451 & ~n_3452;
assign n_3454 =  x_1805 & ~n_3453;
assign n_3455 = ~x_1805 &  n_3453;
assign n_3456 = ~n_3454 & ~n_3455;
assign n_3457 =  x_1804 & ~n_3276;
assign n_3458 =  i_2 &  n_3276;
assign n_3459 = ~n_3457 & ~n_3458;
assign n_3460 =  x_1804 & ~n_3459;
assign n_3461 = ~x_1804 &  n_3459;
assign n_3462 = ~n_3460 & ~n_3461;
assign n_3463 =  x_1803 & ~n_3276;
assign n_3464 =  i_1 &  n_3276;
assign n_3465 = ~n_3463 & ~n_3464;
assign n_3466 =  x_1803 & ~n_3465;
assign n_3467 = ~x_1803 &  n_3465;
assign n_3468 = ~n_3466 & ~n_3467;
assign n_3469 =  x_41 &  n_386;
assign n_3470 =  n_3469 &  n_588;
assign n_3471 =  x_1802 & ~n_3470;
assign n_3472 =  i_32 &  n_3470;
assign n_3473 = ~n_3471 & ~n_3472;
assign n_3474 =  x_1802 & ~n_3473;
assign n_3475 = ~x_1802 &  n_3473;
assign n_3476 = ~n_3474 & ~n_3475;
assign n_3477 =  x_1801 & ~n_3470;
assign n_3478 =  i_31 &  n_3470;
assign n_3479 = ~n_3477 & ~n_3478;
assign n_3480 =  x_1801 & ~n_3479;
assign n_3481 = ~x_1801 &  n_3479;
assign n_3482 = ~n_3480 & ~n_3481;
assign n_3483 =  x_1800 & ~n_3470;
assign n_3484 =  i_30 &  n_3470;
assign n_3485 = ~n_3483 & ~n_3484;
assign n_3486 =  x_1800 & ~n_3485;
assign n_3487 = ~x_1800 &  n_3485;
assign n_3488 = ~n_3486 & ~n_3487;
assign n_3489 =  x_1799 & ~n_3470;
assign n_3490 =  i_29 &  n_3470;
assign n_3491 = ~n_3489 & ~n_3490;
assign n_3492 =  x_1799 & ~n_3491;
assign n_3493 = ~x_1799 &  n_3491;
assign n_3494 = ~n_3492 & ~n_3493;
assign n_3495 =  x_1798 & ~n_3470;
assign n_3496 =  i_28 &  n_3470;
assign n_3497 = ~n_3495 & ~n_3496;
assign n_3498 =  x_1798 & ~n_3497;
assign n_3499 = ~x_1798 &  n_3497;
assign n_3500 = ~n_3498 & ~n_3499;
assign n_3501 =  x_1797 & ~n_3470;
assign n_3502 =  i_27 &  n_3470;
assign n_3503 = ~n_3501 & ~n_3502;
assign n_3504 =  x_1797 & ~n_3503;
assign n_3505 = ~x_1797 &  n_3503;
assign n_3506 = ~n_3504 & ~n_3505;
assign n_3507 =  x_1796 & ~n_3470;
assign n_3508 =  i_26 &  n_3470;
assign n_3509 = ~n_3507 & ~n_3508;
assign n_3510 =  x_1796 & ~n_3509;
assign n_3511 = ~x_1796 &  n_3509;
assign n_3512 = ~n_3510 & ~n_3511;
assign n_3513 =  x_1795 & ~n_3470;
assign n_3514 =  i_25 &  n_3470;
assign n_3515 = ~n_3513 & ~n_3514;
assign n_3516 =  x_1795 & ~n_3515;
assign n_3517 = ~x_1795 &  n_3515;
assign n_3518 = ~n_3516 & ~n_3517;
assign n_3519 =  x_1794 & ~n_3470;
assign n_3520 =  i_24 &  n_3470;
assign n_3521 = ~n_3519 & ~n_3520;
assign n_3522 =  x_1794 & ~n_3521;
assign n_3523 = ~x_1794 &  n_3521;
assign n_3524 = ~n_3522 & ~n_3523;
assign n_3525 =  x_1793 & ~n_3470;
assign n_3526 =  i_23 &  n_3470;
assign n_3527 = ~n_3525 & ~n_3526;
assign n_3528 =  x_1793 & ~n_3527;
assign n_3529 = ~x_1793 &  n_3527;
assign n_3530 = ~n_3528 & ~n_3529;
assign n_3531 =  x_1792 & ~n_3470;
assign n_3532 =  i_22 &  n_3470;
assign n_3533 = ~n_3531 & ~n_3532;
assign n_3534 =  x_1792 & ~n_3533;
assign n_3535 = ~x_1792 &  n_3533;
assign n_3536 = ~n_3534 & ~n_3535;
assign n_3537 =  x_1791 & ~n_3470;
assign n_3538 =  i_21 &  n_3470;
assign n_3539 = ~n_3537 & ~n_3538;
assign n_3540 =  x_1791 & ~n_3539;
assign n_3541 = ~x_1791 &  n_3539;
assign n_3542 = ~n_3540 & ~n_3541;
assign n_3543 =  x_1790 & ~n_3470;
assign n_3544 =  i_20 &  n_3470;
assign n_3545 = ~n_3543 & ~n_3544;
assign n_3546 =  x_1790 & ~n_3545;
assign n_3547 = ~x_1790 &  n_3545;
assign n_3548 = ~n_3546 & ~n_3547;
assign n_3549 =  x_1789 & ~n_3470;
assign n_3550 =  i_19 &  n_3470;
assign n_3551 = ~n_3549 & ~n_3550;
assign n_3552 =  x_1789 & ~n_3551;
assign n_3553 = ~x_1789 &  n_3551;
assign n_3554 = ~n_3552 & ~n_3553;
assign n_3555 =  x_1788 & ~n_3470;
assign n_3556 =  i_18 &  n_3470;
assign n_3557 = ~n_3555 & ~n_3556;
assign n_3558 =  x_1788 & ~n_3557;
assign n_3559 = ~x_1788 &  n_3557;
assign n_3560 = ~n_3558 & ~n_3559;
assign n_3561 =  x_1787 & ~n_3470;
assign n_3562 =  i_17 &  n_3470;
assign n_3563 = ~n_3561 & ~n_3562;
assign n_3564 =  x_1787 & ~n_3563;
assign n_3565 = ~x_1787 &  n_3563;
assign n_3566 = ~n_3564 & ~n_3565;
assign n_3567 =  x_1786 & ~n_3470;
assign n_3568 =  i_16 &  n_3470;
assign n_3569 = ~n_3567 & ~n_3568;
assign n_3570 =  x_1786 & ~n_3569;
assign n_3571 = ~x_1786 &  n_3569;
assign n_3572 = ~n_3570 & ~n_3571;
assign n_3573 =  x_1785 & ~n_3470;
assign n_3574 =  i_15 &  n_3470;
assign n_3575 = ~n_3573 & ~n_3574;
assign n_3576 =  x_1785 & ~n_3575;
assign n_3577 = ~x_1785 &  n_3575;
assign n_3578 = ~n_3576 & ~n_3577;
assign n_3579 =  x_1784 & ~n_3470;
assign n_3580 =  i_14 &  n_3470;
assign n_3581 = ~n_3579 & ~n_3580;
assign n_3582 =  x_1784 & ~n_3581;
assign n_3583 = ~x_1784 &  n_3581;
assign n_3584 = ~n_3582 & ~n_3583;
assign n_3585 =  x_1783 & ~n_3470;
assign n_3586 =  i_13 &  n_3470;
assign n_3587 = ~n_3585 & ~n_3586;
assign n_3588 =  x_1783 & ~n_3587;
assign n_3589 = ~x_1783 &  n_3587;
assign n_3590 = ~n_3588 & ~n_3589;
assign n_3591 =  x_1782 & ~n_3470;
assign n_3592 =  i_12 &  n_3470;
assign n_3593 = ~n_3591 & ~n_3592;
assign n_3594 =  x_1782 & ~n_3593;
assign n_3595 = ~x_1782 &  n_3593;
assign n_3596 = ~n_3594 & ~n_3595;
assign n_3597 =  x_1781 & ~n_3470;
assign n_3598 =  i_11 &  n_3470;
assign n_3599 = ~n_3597 & ~n_3598;
assign n_3600 =  x_1781 & ~n_3599;
assign n_3601 = ~x_1781 &  n_3599;
assign n_3602 = ~n_3600 & ~n_3601;
assign n_3603 =  x_1780 & ~n_3470;
assign n_3604 =  i_10 &  n_3470;
assign n_3605 = ~n_3603 & ~n_3604;
assign n_3606 =  x_1780 & ~n_3605;
assign n_3607 = ~x_1780 &  n_3605;
assign n_3608 = ~n_3606 & ~n_3607;
assign n_3609 =  x_1779 & ~n_3470;
assign n_3610 =  i_9 &  n_3470;
assign n_3611 = ~n_3609 & ~n_3610;
assign n_3612 =  x_1779 & ~n_3611;
assign n_3613 = ~x_1779 &  n_3611;
assign n_3614 = ~n_3612 & ~n_3613;
assign n_3615 =  x_1778 & ~n_3470;
assign n_3616 =  i_8 &  n_3470;
assign n_3617 = ~n_3615 & ~n_3616;
assign n_3618 =  x_1778 & ~n_3617;
assign n_3619 = ~x_1778 &  n_3617;
assign n_3620 = ~n_3618 & ~n_3619;
assign n_3621 =  x_1777 & ~n_3470;
assign n_3622 =  i_7 &  n_3470;
assign n_3623 = ~n_3621 & ~n_3622;
assign n_3624 =  x_1777 & ~n_3623;
assign n_3625 = ~x_1777 &  n_3623;
assign n_3626 = ~n_3624 & ~n_3625;
assign n_3627 =  x_1776 & ~n_3470;
assign n_3628 =  i_6 &  n_3470;
assign n_3629 = ~n_3627 & ~n_3628;
assign n_3630 =  x_1776 & ~n_3629;
assign n_3631 = ~x_1776 &  n_3629;
assign n_3632 = ~n_3630 & ~n_3631;
assign n_3633 =  x_1775 & ~n_3470;
assign n_3634 =  i_5 &  n_3470;
assign n_3635 = ~n_3633 & ~n_3634;
assign n_3636 =  x_1775 & ~n_3635;
assign n_3637 = ~x_1775 &  n_3635;
assign n_3638 = ~n_3636 & ~n_3637;
assign n_3639 =  x_1774 & ~n_3470;
assign n_3640 =  i_4 &  n_3470;
assign n_3641 = ~n_3639 & ~n_3640;
assign n_3642 =  x_1774 & ~n_3641;
assign n_3643 = ~x_1774 &  n_3641;
assign n_3644 = ~n_3642 & ~n_3643;
assign n_3645 =  x_1773 & ~n_3470;
assign n_3646 =  i_3 &  n_3470;
assign n_3647 = ~n_3645 & ~n_3646;
assign n_3648 =  x_1773 & ~n_3647;
assign n_3649 = ~x_1773 &  n_3647;
assign n_3650 = ~n_3648 & ~n_3649;
assign n_3651 =  x_1772 & ~n_3470;
assign n_3652 =  i_2 &  n_3470;
assign n_3653 = ~n_3651 & ~n_3652;
assign n_3654 =  x_1772 & ~n_3653;
assign n_3655 = ~x_1772 &  n_3653;
assign n_3656 = ~n_3654 & ~n_3655;
assign n_3657 =  x_1771 & ~n_3470;
assign n_3658 =  i_1 &  n_3470;
assign n_3659 = ~n_3657 & ~n_3658;
assign n_3660 =  x_1771 & ~n_3659;
assign n_3661 = ~x_1771 &  n_3659;
assign n_3662 = ~n_3660 & ~n_3661;
assign n_3663 = ~x_41 &  n_385;
assign n_3664 =  x_42 &  n_3663;
assign n_3665 =  n_3664 &  n_588;
assign n_3666 =  x_1770 & ~n_3665;
assign n_3667 =  i_32 &  n_3665;
assign n_3668 = ~n_3666 & ~n_3667;
assign n_3669 =  x_1770 & ~n_3668;
assign n_3670 = ~x_1770 &  n_3668;
assign n_3671 = ~n_3669 & ~n_3670;
assign n_3672 =  x_1769 & ~n_3665;
assign n_3673 =  i_31 &  n_3665;
assign n_3674 = ~n_3672 & ~n_3673;
assign n_3675 =  x_1769 & ~n_3674;
assign n_3676 = ~x_1769 &  n_3674;
assign n_3677 = ~n_3675 & ~n_3676;
assign n_3678 =  x_1768 & ~n_3665;
assign n_3679 =  i_30 &  n_3665;
assign n_3680 = ~n_3678 & ~n_3679;
assign n_3681 =  x_1768 & ~n_3680;
assign n_3682 = ~x_1768 &  n_3680;
assign n_3683 = ~n_3681 & ~n_3682;
assign n_3684 =  x_1767 & ~n_3665;
assign n_3685 =  i_29 &  n_3665;
assign n_3686 = ~n_3684 & ~n_3685;
assign n_3687 =  x_1767 & ~n_3686;
assign n_3688 = ~x_1767 &  n_3686;
assign n_3689 = ~n_3687 & ~n_3688;
assign n_3690 =  x_1766 & ~n_3665;
assign n_3691 =  i_28 &  n_3665;
assign n_3692 = ~n_3690 & ~n_3691;
assign n_3693 =  x_1766 & ~n_3692;
assign n_3694 = ~x_1766 &  n_3692;
assign n_3695 = ~n_3693 & ~n_3694;
assign n_3696 =  x_1765 & ~n_3665;
assign n_3697 =  i_27 &  n_3665;
assign n_3698 = ~n_3696 & ~n_3697;
assign n_3699 =  x_1765 & ~n_3698;
assign n_3700 = ~x_1765 &  n_3698;
assign n_3701 = ~n_3699 & ~n_3700;
assign n_3702 =  x_1764 & ~n_3665;
assign n_3703 =  i_26 &  n_3665;
assign n_3704 = ~n_3702 & ~n_3703;
assign n_3705 =  x_1764 & ~n_3704;
assign n_3706 = ~x_1764 &  n_3704;
assign n_3707 = ~n_3705 & ~n_3706;
assign n_3708 =  x_1763 & ~n_3665;
assign n_3709 =  i_25 &  n_3665;
assign n_3710 = ~n_3708 & ~n_3709;
assign n_3711 =  x_1763 & ~n_3710;
assign n_3712 = ~x_1763 &  n_3710;
assign n_3713 = ~n_3711 & ~n_3712;
assign n_3714 =  x_1762 & ~n_3665;
assign n_3715 =  i_24 &  n_3665;
assign n_3716 = ~n_3714 & ~n_3715;
assign n_3717 =  x_1762 & ~n_3716;
assign n_3718 = ~x_1762 &  n_3716;
assign n_3719 = ~n_3717 & ~n_3718;
assign n_3720 =  x_1761 & ~n_3665;
assign n_3721 =  i_23 &  n_3665;
assign n_3722 = ~n_3720 & ~n_3721;
assign n_3723 =  x_1761 & ~n_3722;
assign n_3724 = ~x_1761 &  n_3722;
assign n_3725 = ~n_3723 & ~n_3724;
assign n_3726 =  x_1760 & ~n_3665;
assign n_3727 =  i_22 &  n_3665;
assign n_3728 = ~n_3726 & ~n_3727;
assign n_3729 =  x_1760 & ~n_3728;
assign n_3730 = ~x_1760 &  n_3728;
assign n_3731 = ~n_3729 & ~n_3730;
assign n_3732 =  x_1759 & ~n_3665;
assign n_3733 =  i_21 &  n_3665;
assign n_3734 = ~n_3732 & ~n_3733;
assign n_3735 =  x_1759 & ~n_3734;
assign n_3736 = ~x_1759 &  n_3734;
assign n_3737 = ~n_3735 & ~n_3736;
assign n_3738 =  x_1758 & ~n_3665;
assign n_3739 =  i_20 &  n_3665;
assign n_3740 = ~n_3738 & ~n_3739;
assign n_3741 =  x_1758 & ~n_3740;
assign n_3742 = ~x_1758 &  n_3740;
assign n_3743 = ~n_3741 & ~n_3742;
assign n_3744 =  x_1757 & ~n_3665;
assign n_3745 =  i_19 &  n_3665;
assign n_3746 = ~n_3744 & ~n_3745;
assign n_3747 =  x_1757 & ~n_3746;
assign n_3748 = ~x_1757 &  n_3746;
assign n_3749 = ~n_3747 & ~n_3748;
assign n_3750 =  x_1756 & ~n_3665;
assign n_3751 =  i_18 &  n_3665;
assign n_3752 = ~n_3750 & ~n_3751;
assign n_3753 =  x_1756 & ~n_3752;
assign n_3754 = ~x_1756 &  n_3752;
assign n_3755 = ~n_3753 & ~n_3754;
assign n_3756 =  x_1755 & ~n_3665;
assign n_3757 =  i_17 &  n_3665;
assign n_3758 = ~n_3756 & ~n_3757;
assign n_3759 =  x_1755 & ~n_3758;
assign n_3760 = ~x_1755 &  n_3758;
assign n_3761 = ~n_3759 & ~n_3760;
assign n_3762 =  x_1754 & ~n_3665;
assign n_3763 =  i_16 &  n_3665;
assign n_3764 = ~n_3762 & ~n_3763;
assign n_3765 =  x_1754 & ~n_3764;
assign n_3766 = ~x_1754 &  n_3764;
assign n_3767 = ~n_3765 & ~n_3766;
assign n_3768 =  x_1753 & ~n_3665;
assign n_3769 =  i_15 &  n_3665;
assign n_3770 = ~n_3768 & ~n_3769;
assign n_3771 =  x_1753 & ~n_3770;
assign n_3772 = ~x_1753 &  n_3770;
assign n_3773 = ~n_3771 & ~n_3772;
assign n_3774 =  x_1752 & ~n_3665;
assign n_3775 =  i_14 &  n_3665;
assign n_3776 = ~n_3774 & ~n_3775;
assign n_3777 =  x_1752 & ~n_3776;
assign n_3778 = ~x_1752 &  n_3776;
assign n_3779 = ~n_3777 & ~n_3778;
assign n_3780 =  x_1751 & ~n_3665;
assign n_3781 =  i_13 &  n_3665;
assign n_3782 = ~n_3780 & ~n_3781;
assign n_3783 =  x_1751 & ~n_3782;
assign n_3784 = ~x_1751 &  n_3782;
assign n_3785 = ~n_3783 & ~n_3784;
assign n_3786 =  x_1750 & ~n_3665;
assign n_3787 =  i_12 &  n_3665;
assign n_3788 = ~n_3786 & ~n_3787;
assign n_3789 =  x_1750 & ~n_3788;
assign n_3790 = ~x_1750 &  n_3788;
assign n_3791 = ~n_3789 & ~n_3790;
assign n_3792 =  x_1749 & ~n_3665;
assign n_3793 =  i_11 &  n_3665;
assign n_3794 = ~n_3792 & ~n_3793;
assign n_3795 =  x_1749 & ~n_3794;
assign n_3796 = ~x_1749 &  n_3794;
assign n_3797 = ~n_3795 & ~n_3796;
assign n_3798 =  x_1748 & ~n_3665;
assign n_3799 =  i_10 &  n_3665;
assign n_3800 = ~n_3798 & ~n_3799;
assign n_3801 =  x_1748 & ~n_3800;
assign n_3802 = ~x_1748 &  n_3800;
assign n_3803 = ~n_3801 & ~n_3802;
assign n_3804 =  x_1747 & ~n_3665;
assign n_3805 =  i_9 &  n_3665;
assign n_3806 = ~n_3804 & ~n_3805;
assign n_3807 =  x_1747 & ~n_3806;
assign n_3808 = ~x_1747 &  n_3806;
assign n_3809 = ~n_3807 & ~n_3808;
assign n_3810 =  x_1746 & ~n_3665;
assign n_3811 =  i_8 &  n_3665;
assign n_3812 = ~n_3810 & ~n_3811;
assign n_3813 =  x_1746 & ~n_3812;
assign n_3814 = ~x_1746 &  n_3812;
assign n_3815 = ~n_3813 & ~n_3814;
assign n_3816 =  x_1745 & ~n_3665;
assign n_3817 =  i_7 &  n_3665;
assign n_3818 = ~n_3816 & ~n_3817;
assign n_3819 =  x_1745 & ~n_3818;
assign n_3820 = ~x_1745 &  n_3818;
assign n_3821 = ~n_3819 & ~n_3820;
assign n_3822 =  x_1744 & ~n_3665;
assign n_3823 =  i_6 &  n_3665;
assign n_3824 = ~n_3822 & ~n_3823;
assign n_3825 =  x_1744 & ~n_3824;
assign n_3826 = ~x_1744 &  n_3824;
assign n_3827 = ~n_3825 & ~n_3826;
assign n_3828 =  x_1743 & ~n_3665;
assign n_3829 =  i_5 &  n_3665;
assign n_3830 = ~n_3828 & ~n_3829;
assign n_3831 =  x_1743 & ~n_3830;
assign n_3832 = ~x_1743 &  n_3830;
assign n_3833 = ~n_3831 & ~n_3832;
assign n_3834 =  x_1742 & ~n_3665;
assign n_3835 =  i_4 &  n_3665;
assign n_3836 = ~n_3834 & ~n_3835;
assign n_3837 =  x_1742 & ~n_3836;
assign n_3838 = ~x_1742 &  n_3836;
assign n_3839 = ~n_3837 & ~n_3838;
assign n_3840 =  x_1741 & ~n_3665;
assign n_3841 =  i_3 &  n_3665;
assign n_3842 = ~n_3840 & ~n_3841;
assign n_3843 =  x_1741 & ~n_3842;
assign n_3844 = ~x_1741 &  n_3842;
assign n_3845 = ~n_3843 & ~n_3844;
assign n_3846 =  x_1740 & ~n_3665;
assign n_3847 =  i_2 &  n_3665;
assign n_3848 = ~n_3846 & ~n_3847;
assign n_3849 =  x_1740 & ~n_3848;
assign n_3850 = ~x_1740 &  n_3848;
assign n_3851 = ~n_3849 & ~n_3850;
assign n_3852 =  x_1739 & ~n_3665;
assign n_3853 =  i_1 &  n_3665;
assign n_3854 = ~n_3852 & ~n_3853;
assign n_3855 =  x_1739 & ~n_3854;
assign n_3856 = ~x_1739 &  n_3854;
assign n_3857 = ~n_3855 & ~n_3856;
assign n_3858 = ~x_42 &  n_1;
assign n_3859 =  x_36 &  x_37;
assign n_3860 =  n_387 &  n_3859;
assign n_3861 = ~x_38 & ~x_39;
assign n_3862 =  n_3860 &  n_3861;
assign n_3863 =  n_3858 &  n_3862;
assign n_3864 =  x_1738 & ~n_3863;
assign n_3865 =  i_32 &  n_3863;
assign n_3866 = ~n_3864 & ~n_3865;
assign n_3867 =  x_1738 & ~n_3866;
assign n_3868 = ~x_1738 &  n_3866;
assign n_3869 = ~n_3867 & ~n_3868;
assign n_3870 =  x_1737 & ~n_3863;
assign n_3871 =  i_31 &  n_3863;
assign n_3872 = ~n_3870 & ~n_3871;
assign n_3873 =  x_1737 & ~n_3872;
assign n_3874 = ~x_1737 &  n_3872;
assign n_3875 = ~n_3873 & ~n_3874;
assign n_3876 =  x_1736 & ~n_3863;
assign n_3877 =  i_30 &  n_3863;
assign n_3878 = ~n_3876 & ~n_3877;
assign n_3879 =  x_1736 & ~n_3878;
assign n_3880 = ~x_1736 &  n_3878;
assign n_3881 = ~n_3879 & ~n_3880;
assign n_3882 =  x_1735 & ~n_3863;
assign n_3883 =  i_29 &  n_3863;
assign n_3884 = ~n_3882 & ~n_3883;
assign n_3885 =  x_1735 & ~n_3884;
assign n_3886 = ~x_1735 &  n_3884;
assign n_3887 = ~n_3885 & ~n_3886;
assign n_3888 =  x_1734 & ~n_3863;
assign n_3889 =  i_28 &  n_3863;
assign n_3890 = ~n_3888 & ~n_3889;
assign n_3891 =  x_1734 & ~n_3890;
assign n_3892 = ~x_1734 &  n_3890;
assign n_3893 = ~n_3891 & ~n_3892;
assign n_3894 =  x_1733 & ~n_3863;
assign n_3895 =  i_27 &  n_3863;
assign n_3896 = ~n_3894 & ~n_3895;
assign n_3897 =  x_1733 & ~n_3896;
assign n_3898 = ~x_1733 &  n_3896;
assign n_3899 = ~n_3897 & ~n_3898;
assign n_3900 =  x_1732 & ~n_3863;
assign n_3901 =  i_26 &  n_3863;
assign n_3902 = ~n_3900 & ~n_3901;
assign n_3903 =  x_1732 & ~n_3902;
assign n_3904 = ~x_1732 &  n_3902;
assign n_3905 = ~n_3903 & ~n_3904;
assign n_3906 =  x_1731 & ~n_3863;
assign n_3907 =  i_25 &  n_3863;
assign n_3908 = ~n_3906 & ~n_3907;
assign n_3909 =  x_1731 & ~n_3908;
assign n_3910 = ~x_1731 &  n_3908;
assign n_3911 = ~n_3909 & ~n_3910;
assign n_3912 =  x_1730 & ~n_3863;
assign n_3913 =  i_24 &  n_3863;
assign n_3914 = ~n_3912 & ~n_3913;
assign n_3915 =  x_1730 & ~n_3914;
assign n_3916 = ~x_1730 &  n_3914;
assign n_3917 = ~n_3915 & ~n_3916;
assign n_3918 =  x_1729 & ~n_3863;
assign n_3919 =  i_23 &  n_3863;
assign n_3920 = ~n_3918 & ~n_3919;
assign n_3921 =  x_1729 & ~n_3920;
assign n_3922 = ~x_1729 &  n_3920;
assign n_3923 = ~n_3921 & ~n_3922;
assign n_3924 =  x_1728 & ~n_3863;
assign n_3925 =  i_22 &  n_3863;
assign n_3926 = ~n_3924 & ~n_3925;
assign n_3927 =  x_1728 & ~n_3926;
assign n_3928 = ~x_1728 &  n_3926;
assign n_3929 = ~n_3927 & ~n_3928;
assign n_3930 =  x_1727 & ~n_3863;
assign n_3931 =  i_21 &  n_3863;
assign n_3932 = ~n_3930 & ~n_3931;
assign n_3933 =  x_1727 & ~n_3932;
assign n_3934 = ~x_1727 &  n_3932;
assign n_3935 = ~n_3933 & ~n_3934;
assign n_3936 =  x_1726 & ~n_3863;
assign n_3937 =  i_20 &  n_3863;
assign n_3938 = ~n_3936 & ~n_3937;
assign n_3939 =  x_1726 & ~n_3938;
assign n_3940 = ~x_1726 &  n_3938;
assign n_3941 = ~n_3939 & ~n_3940;
assign n_3942 =  x_1725 & ~n_3863;
assign n_3943 =  i_19 &  n_3863;
assign n_3944 = ~n_3942 & ~n_3943;
assign n_3945 =  x_1725 & ~n_3944;
assign n_3946 = ~x_1725 &  n_3944;
assign n_3947 = ~n_3945 & ~n_3946;
assign n_3948 =  x_1724 & ~n_3863;
assign n_3949 =  i_18 &  n_3863;
assign n_3950 = ~n_3948 & ~n_3949;
assign n_3951 =  x_1724 & ~n_3950;
assign n_3952 = ~x_1724 &  n_3950;
assign n_3953 = ~n_3951 & ~n_3952;
assign n_3954 =  x_1723 & ~n_3863;
assign n_3955 =  i_17 &  n_3863;
assign n_3956 = ~n_3954 & ~n_3955;
assign n_3957 =  x_1723 & ~n_3956;
assign n_3958 = ~x_1723 &  n_3956;
assign n_3959 = ~n_3957 & ~n_3958;
assign n_3960 =  x_1722 & ~n_3863;
assign n_3961 =  i_16 &  n_3863;
assign n_3962 = ~n_3960 & ~n_3961;
assign n_3963 =  x_1722 & ~n_3962;
assign n_3964 = ~x_1722 &  n_3962;
assign n_3965 = ~n_3963 & ~n_3964;
assign n_3966 =  x_1721 & ~n_3863;
assign n_3967 =  i_15 &  n_3863;
assign n_3968 = ~n_3966 & ~n_3967;
assign n_3969 =  x_1721 & ~n_3968;
assign n_3970 = ~x_1721 &  n_3968;
assign n_3971 = ~n_3969 & ~n_3970;
assign n_3972 =  x_1720 & ~n_3863;
assign n_3973 =  i_14 &  n_3863;
assign n_3974 = ~n_3972 & ~n_3973;
assign n_3975 =  x_1720 & ~n_3974;
assign n_3976 = ~x_1720 &  n_3974;
assign n_3977 = ~n_3975 & ~n_3976;
assign n_3978 =  x_1719 & ~n_3863;
assign n_3979 =  i_13 &  n_3863;
assign n_3980 = ~n_3978 & ~n_3979;
assign n_3981 =  x_1719 & ~n_3980;
assign n_3982 = ~x_1719 &  n_3980;
assign n_3983 = ~n_3981 & ~n_3982;
assign n_3984 =  x_1718 & ~n_3863;
assign n_3985 =  i_12 &  n_3863;
assign n_3986 = ~n_3984 & ~n_3985;
assign n_3987 =  x_1718 & ~n_3986;
assign n_3988 = ~x_1718 &  n_3986;
assign n_3989 = ~n_3987 & ~n_3988;
assign n_3990 =  x_1717 & ~n_3863;
assign n_3991 =  i_11 &  n_3863;
assign n_3992 = ~n_3990 & ~n_3991;
assign n_3993 =  x_1717 & ~n_3992;
assign n_3994 = ~x_1717 &  n_3992;
assign n_3995 = ~n_3993 & ~n_3994;
assign n_3996 =  x_1716 & ~n_3863;
assign n_3997 =  i_10 &  n_3863;
assign n_3998 = ~n_3996 & ~n_3997;
assign n_3999 =  x_1716 & ~n_3998;
assign n_4000 = ~x_1716 &  n_3998;
assign n_4001 = ~n_3999 & ~n_4000;
assign n_4002 =  x_1715 & ~n_3863;
assign n_4003 =  i_9 &  n_3863;
assign n_4004 = ~n_4002 & ~n_4003;
assign n_4005 =  x_1715 & ~n_4004;
assign n_4006 = ~x_1715 &  n_4004;
assign n_4007 = ~n_4005 & ~n_4006;
assign n_4008 =  x_1714 & ~n_3863;
assign n_4009 =  i_8 &  n_3863;
assign n_4010 = ~n_4008 & ~n_4009;
assign n_4011 =  x_1714 & ~n_4010;
assign n_4012 = ~x_1714 &  n_4010;
assign n_4013 = ~n_4011 & ~n_4012;
assign n_4014 =  x_1713 & ~n_3863;
assign n_4015 =  i_7 &  n_3863;
assign n_4016 = ~n_4014 & ~n_4015;
assign n_4017 =  x_1713 & ~n_4016;
assign n_4018 = ~x_1713 &  n_4016;
assign n_4019 = ~n_4017 & ~n_4018;
assign n_4020 =  x_1712 & ~n_3863;
assign n_4021 =  i_6 &  n_3863;
assign n_4022 = ~n_4020 & ~n_4021;
assign n_4023 =  x_1712 & ~n_4022;
assign n_4024 = ~x_1712 &  n_4022;
assign n_4025 = ~n_4023 & ~n_4024;
assign n_4026 =  x_1711 & ~n_3863;
assign n_4027 =  i_5 &  n_3863;
assign n_4028 = ~n_4026 & ~n_4027;
assign n_4029 =  x_1711 & ~n_4028;
assign n_4030 = ~x_1711 &  n_4028;
assign n_4031 = ~n_4029 & ~n_4030;
assign n_4032 =  x_1710 & ~n_3863;
assign n_4033 =  i_4 &  n_3863;
assign n_4034 = ~n_4032 & ~n_4033;
assign n_4035 =  x_1710 & ~n_4034;
assign n_4036 = ~x_1710 &  n_4034;
assign n_4037 = ~n_4035 & ~n_4036;
assign n_4038 =  x_1709 & ~n_3863;
assign n_4039 =  i_3 &  n_3863;
assign n_4040 = ~n_4038 & ~n_4039;
assign n_4041 =  x_1709 & ~n_4040;
assign n_4042 = ~x_1709 &  n_4040;
assign n_4043 = ~n_4041 & ~n_4042;
assign n_4044 =  x_1708 & ~n_3863;
assign n_4045 =  i_2 &  n_3863;
assign n_4046 = ~n_4044 & ~n_4045;
assign n_4047 =  x_1708 & ~n_4046;
assign n_4048 = ~x_1708 &  n_4046;
assign n_4049 = ~n_4047 & ~n_4048;
assign n_4050 =  x_1707 & ~n_3863;
assign n_4051 =  i_1 &  n_3863;
assign n_4052 = ~n_4050 & ~n_4051;
assign n_4053 =  x_1707 & ~n_4052;
assign n_4054 = ~x_1707 &  n_4052;
assign n_4055 = ~n_4053 & ~n_4054;
assign n_4056 =  n_188 &  n_389;
assign n_4057 =  n_189 &  n_4056;
assign n_4058 =  n_1707 &  n_4057;
assign n_4059 =  x_1706 & ~n_4058;
assign n_4060 =  i_32 &  n_4058;
assign n_4061 = ~n_4059 & ~n_4060;
assign n_4062 =  x_1706 & ~n_4061;
assign n_4063 = ~x_1706 &  n_4061;
assign n_4064 = ~n_4062 & ~n_4063;
assign n_4065 =  x_1705 & ~n_4058;
assign n_4066 =  i_31 &  n_4058;
assign n_4067 = ~n_4065 & ~n_4066;
assign n_4068 =  x_1705 & ~n_4067;
assign n_4069 = ~x_1705 &  n_4067;
assign n_4070 = ~n_4068 & ~n_4069;
assign n_4071 =  x_1704 & ~n_4058;
assign n_4072 =  i_30 &  n_4058;
assign n_4073 = ~n_4071 & ~n_4072;
assign n_4074 =  x_1704 & ~n_4073;
assign n_4075 = ~x_1704 &  n_4073;
assign n_4076 = ~n_4074 & ~n_4075;
assign n_4077 =  x_1703 & ~n_4058;
assign n_4078 =  i_29 &  n_4058;
assign n_4079 = ~n_4077 & ~n_4078;
assign n_4080 =  x_1703 & ~n_4079;
assign n_4081 = ~x_1703 &  n_4079;
assign n_4082 = ~n_4080 & ~n_4081;
assign n_4083 =  x_1702 & ~n_4058;
assign n_4084 =  i_28 &  n_4058;
assign n_4085 = ~n_4083 & ~n_4084;
assign n_4086 =  x_1702 & ~n_4085;
assign n_4087 = ~x_1702 &  n_4085;
assign n_4088 = ~n_4086 & ~n_4087;
assign n_4089 =  x_1701 & ~n_4058;
assign n_4090 =  i_27 &  n_4058;
assign n_4091 = ~n_4089 & ~n_4090;
assign n_4092 =  x_1701 & ~n_4091;
assign n_4093 = ~x_1701 &  n_4091;
assign n_4094 = ~n_4092 & ~n_4093;
assign n_4095 =  x_1700 & ~n_4058;
assign n_4096 =  i_26 &  n_4058;
assign n_4097 = ~n_4095 & ~n_4096;
assign n_4098 =  x_1700 & ~n_4097;
assign n_4099 = ~x_1700 &  n_4097;
assign n_4100 = ~n_4098 & ~n_4099;
assign n_4101 =  x_1699 & ~n_4058;
assign n_4102 =  i_25 &  n_4058;
assign n_4103 = ~n_4101 & ~n_4102;
assign n_4104 =  x_1699 & ~n_4103;
assign n_4105 = ~x_1699 &  n_4103;
assign n_4106 = ~n_4104 & ~n_4105;
assign n_4107 =  x_1698 & ~n_4058;
assign n_4108 =  i_24 &  n_4058;
assign n_4109 = ~n_4107 & ~n_4108;
assign n_4110 =  x_1698 & ~n_4109;
assign n_4111 = ~x_1698 &  n_4109;
assign n_4112 = ~n_4110 & ~n_4111;
assign n_4113 =  x_1697 & ~n_4058;
assign n_4114 =  i_23 &  n_4058;
assign n_4115 = ~n_4113 & ~n_4114;
assign n_4116 =  x_1697 & ~n_4115;
assign n_4117 = ~x_1697 &  n_4115;
assign n_4118 = ~n_4116 & ~n_4117;
assign n_4119 =  x_1696 & ~n_4058;
assign n_4120 =  i_22 &  n_4058;
assign n_4121 = ~n_4119 & ~n_4120;
assign n_4122 =  x_1696 & ~n_4121;
assign n_4123 = ~x_1696 &  n_4121;
assign n_4124 = ~n_4122 & ~n_4123;
assign n_4125 =  x_1695 & ~n_4058;
assign n_4126 =  i_21 &  n_4058;
assign n_4127 = ~n_4125 & ~n_4126;
assign n_4128 =  x_1695 & ~n_4127;
assign n_4129 = ~x_1695 &  n_4127;
assign n_4130 = ~n_4128 & ~n_4129;
assign n_4131 =  x_1694 & ~n_4058;
assign n_4132 =  i_20 &  n_4058;
assign n_4133 = ~n_4131 & ~n_4132;
assign n_4134 =  x_1694 & ~n_4133;
assign n_4135 = ~x_1694 &  n_4133;
assign n_4136 = ~n_4134 & ~n_4135;
assign n_4137 =  x_1693 & ~n_4058;
assign n_4138 =  i_19 &  n_4058;
assign n_4139 = ~n_4137 & ~n_4138;
assign n_4140 =  x_1693 & ~n_4139;
assign n_4141 = ~x_1693 &  n_4139;
assign n_4142 = ~n_4140 & ~n_4141;
assign n_4143 =  x_1692 & ~n_4058;
assign n_4144 =  i_18 &  n_4058;
assign n_4145 = ~n_4143 & ~n_4144;
assign n_4146 =  x_1692 & ~n_4145;
assign n_4147 = ~x_1692 &  n_4145;
assign n_4148 = ~n_4146 & ~n_4147;
assign n_4149 =  x_1691 & ~n_4058;
assign n_4150 =  i_17 &  n_4058;
assign n_4151 = ~n_4149 & ~n_4150;
assign n_4152 =  x_1691 & ~n_4151;
assign n_4153 = ~x_1691 &  n_4151;
assign n_4154 = ~n_4152 & ~n_4153;
assign n_4155 =  x_1690 & ~n_4058;
assign n_4156 =  i_16 &  n_4058;
assign n_4157 = ~n_4155 & ~n_4156;
assign n_4158 =  x_1690 & ~n_4157;
assign n_4159 = ~x_1690 &  n_4157;
assign n_4160 = ~n_4158 & ~n_4159;
assign n_4161 =  x_1689 & ~n_4058;
assign n_4162 =  i_15 &  n_4058;
assign n_4163 = ~n_4161 & ~n_4162;
assign n_4164 =  x_1689 & ~n_4163;
assign n_4165 = ~x_1689 &  n_4163;
assign n_4166 = ~n_4164 & ~n_4165;
assign n_4167 =  x_1688 & ~n_4058;
assign n_4168 =  i_14 &  n_4058;
assign n_4169 = ~n_4167 & ~n_4168;
assign n_4170 =  x_1688 & ~n_4169;
assign n_4171 = ~x_1688 &  n_4169;
assign n_4172 = ~n_4170 & ~n_4171;
assign n_4173 =  x_1687 & ~n_4058;
assign n_4174 =  i_13 &  n_4058;
assign n_4175 = ~n_4173 & ~n_4174;
assign n_4176 =  x_1687 & ~n_4175;
assign n_4177 = ~x_1687 &  n_4175;
assign n_4178 = ~n_4176 & ~n_4177;
assign n_4179 =  x_1686 & ~n_4058;
assign n_4180 =  i_12 &  n_4058;
assign n_4181 = ~n_4179 & ~n_4180;
assign n_4182 =  x_1686 & ~n_4181;
assign n_4183 = ~x_1686 &  n_4181;
assign n_4184 = ~n_4182 & ~n_4183;
assign n_4185 =  x_1685 & ~n_4058;
assign n_4186 =  i_11 &  n_4058;
assign n_4187 = ~n_4185 & ~n_4186;
assign n_4188 =  x_1685 & ~n_4187;
assign n_4189 = ~x_1685 &  n_4187;
assign n_4190 = ~n_4188 & ~n_4189;
assign n_4191 =  x_1684 & ~n_4058;
assign n_4192 =  i_10 &  n_4058;
assign n_4193 = ~n_4191 & ~n_4192;
assign n_4194 =  x_1684 & ~n_4193;
assign n_4195 = ~x_1684 &  n_4193;
assign n_4196 = ~n_4194 & ~n_4195;
assign n_4197 =  x_1683 & ~n_4058;
assign n_4198 =  i_9 &  n_4058;
assign n_4199 = ~n_4197 & ~n_4198;
assign n_4200 =  x_1683 & ~n_4199;
assign n_4201 = ~x_1683 &  n_4199;
assign n_4202 = ~n_4200 & ~n_4201;
assign n_4203 =  x_1682 & ~n_4058;
assign n_4204 =  i_8 &  n_4058;
assign n_4205 = ~n_4203 & ~n_4204;
assign n_4206 =  x_1682 & ~n_4205;
assign n_4207 = ~x_1682 &  n_4205;
assign n_4208 = ~n_4206 & ~n_4207;
assign n_4209 =  x_1681 & ~n_4058;
assign n_4210 =  i_7 &  n_4058;
assign n_4211 = ~n_4209 & ~n_4210;
assign n_4212 =  x_1681 & ~n_4211;
assign n_4213 = ~x_1681 &  n_4211;
assign n_4214 = ~n_4212 & ~n_4213;
assign n_4215 =  x_1680 & ~n_4058;
assign n_4216 =  i_6 &  n_4058;
assign n_4217 = ~n_4215 & ~n_4216;
assign n_4218 =  x_1680 & ~n_4217;
assign n_4219 = ~x_1680 &  n_4217;
assign n_4220 = ~n_4218 & ~n_4219;
assign n_4221 =  x_1679 & ~n_4058;
assign n_4222 =  i_5 &  n_4058;
assign n_4223 = ~n_4221 & ~n_4222;
assign n_4224 =  x_1679 & ~n_4223;
assign n_4225 = ~x_1679 &  n_4223;
assign n_4226 = ~n_4224 & ~n_4225;
assign n_4227 =  x_1678 & ~n_4058;
assign n_4228 =  i_4 &  n_4058;
assign n_4229 = ~n_4227 & ~n_4228;
assign n_4230 =  x_1678 & ~n_4229;
assign n_4231 = ~x_1678 &  n_4229;
assign n_4232 = ~n_4230 & ~n_4231;
assign n_4233 =  x_1677 & ~n_4058;
assign n_4234 =  i_3 &  n_4058;
assign n_4235 = ~n_4233 & ~n_4234;
assign n_4236 =  x_1677 & ~n_4235;
assign n_4237 = ~x_1677 &  n_4235;
assign n_4238 = ~n_4236 & ~n_4237;
assign n_4239 =  x_1676 & ~n_4058;
assign n_4240 =  i_2 &  n_4058;
assign n_4241 = ~n_4239 & ~n_4240;
assign n_4242 =  x_1676 & ~n_4241;
assign n_4243 = ~x_1676 &  n_4241;
assign n_4244 = ~n_4242 & ~n_4243;
assign n_4245 =  x_1675 & ~n_4058;
assign n_4246 =  i_1 &  n_4058;
assign n_4247 = ~n_4245 & ~n_4246;
assign n_4248 =  x_1675 & ~n_4247;
assign n_4249 = ~x_1675 &  n_4247;
assign n_4250 = ~n_4248 & ~n_4249;
assign n_4251 =  n_1903 &  n_2302;
assign n_4252 =  n_586 &  n_4251;
assign n_4253 =  x_1674 & ~n_4252;
assign n_4254 =  i_32 &  n_4252;
assign n_4255 = ~n_4253 & ~n_4254;
assign n_4256 =  x_1674 & ~n_4255;
assign n_4257 = ~x_1674 &  n_4255;
assign n_4258 = ~n_4256 & ~n_4257;
assign n_4259 =  x_1673 & ~n_4252;
assign n_4260 =  i_31 &  n_4252;
assign n_4261 = ~n_4259 & ~n_4260;
assign n_4262 =  x_1673 & ~n_4261;
assign n_4263 = ~x_1673 &  n_4261;
assign n_4264 = ~n_4262 & ~n_4263;
assign n_4265 =  x_1672 & ~n_4252;
assign n_4266 =  i_30 &  n_4252;
assign n_4267 = ~n_4265 & ~n_4266;
assign n_4268 =  x_1672 & ~n_4267;
assign n_4269 = ~x_1672 &  n_4267;
assign n_4270 = ~n_4268 & ~n_4269;
assign n_4271 =  x_1671 & ~n_4252;
assign n_4272 =  i_29 &  n_4252;
assign n_4273 = ~n_4271 & ~n_4272;
assign n_4274 =  x_1671 & ~n_4273;
assign n_4275 = ~x_1671 &  n_4273;
assign n_4276 = ~n_4274 & ~n_4275;
assign n_4277 =  x_1670 & ~n_4252;
assign n_4278 =  i_28 &  n_4252;
assign n_4279 = ~n_4277 & ~n_4278;
assign n_4280 =  x_1670 & ~n_4279;
assign n_4281 = ~x_1670 &  n_4279;
assign n_4282 = ~n_4280 & ~n_4281;
assign n_4283 =  x_1669 & ~n_4252;
assign n_4284 =  i_27 &  n_4252;
assign n_4285 = ~n_4283 & ~n_4284;
assign n_4286 =  x_1669 & ~n_4285;
assign n_4287 = ~x_1669 &  n_4285;
assign n_4288 = ~n_4286 & ~n_4287;
assign n_4289 =  x_1668 & ~n_4252;
assign n_4290 =  i_26 &  n_4252;
assign n_4291 = ~n_4289 & ~n_4290;
assign n_4292 =  x_1668 & ~n_4291;
assign n_4293 = ~x_1668 &  n_4291;
assign n_4294 = ~n_4292 & ~n_4293;
assign n_4295 =  x_1667 & ~n_4252;
assign n_4296 =  i_25 &  n_4252;
assign n_4297 = ~n_4295 & ~n_4296;
assign n_4298 =  x_1667 & ~n_4297;
assign n_4299 = ~x_1667 &  n_4297;
assign n_4300 = ~n_4298 & ~n_4299;
assign n_4301 =  x_1666 & ~n_4252;
assign n_4302 =  i_24 &  n_4252;
assign n_4303 = ~n_4301 & ~n_4302;
assign n_4304 =  x_1666 & ~n_4303;
assign n_4305 = ~x_1666 &  n_4303;
assign n_4306 = ~n_4304 & ~n_4305;
assign n_4307 =  x_1665 & ~n_4252;
assign n_4308 =  i_23 &  n_4252;
assign n_4309 = ~n_4307 & ~n_4308;
assign n_4310 =  x_1665 & ~n_4309;
assign n_4311 = ~x_1665 &  n_4309;
assign n_4312 = ~n_4310 & ~n_4311;
assign n_4313 =  x_1664 & ~n_4252;
assign n_4314 =  i_22 &  n_4252;
assign n_4315 = ~n_4313 & ~n_4314;
assign n_4316 =  x_1664 & ~n_4315;
assign n_4317 = ~x_1664 &  n_4315;
assign n_4318 = ~n_4316 & ~n_4317;
assign n_4319 =  x_1663 & ~n_4252;
assign n_4320 =  i_21 &  n_4252;
assign n_4321 = ~n_4319 & ~n_4320;
assign n_4322 =  x_1663 & ~n_4321;
assign n_4323 = ~x_1663 &  n_4321;
assign n_4324 = ~n_4322 & ~n_4323;
assign n_4325 =  x_1662 & ~n_4252;
assign n_4326 =  i_20 &  n_4252;
assign n_4327 = ~n_4325 & ~n_4326;
assign n_4328 =  x_1662 & ~n_4327;
assign n_4329 = ~x_1662 &  n_4327;
assign n_4330 = ~n_4328 & ~n_4329;
assign n_4331 =  x_1661 & ~n_4252;
assign n_4332 =  i_19 &  n_4252;
assign n_4333 = ~n_4331 & ~n_4332;
assign n_4334 =  x_1661 & ~n_4333;
assign n_4335 = ~x_1661 &  n_4333;
assign n_4336 = ~n_4334 & ~n_4335;
assign n_4337 =  x_1660 & ~n_4252;
assign n_4338 =  i_18 &  n_4252;
assign n_4339 = ~n_4337 & ~n_4338;
assign n_4340 =  x_1660 & ~n_4339;
assign n_4341 = ~x_1660 &  n_4339;
assign n_4342 = ~n_4340 & ~n_4341;
assign n_4343 =  x_1659 & ~n_4252;
assign n_4344 =  i_17 &  n_4252;
assign n_4345 = ~n_4343 & ~n_4344;
assign n_4346 =  x_1659 & ~n_4345;
assign n_4347 = ~x_1659 &  n_4345;
assign n_4348 = ~n_4346 & ~n_4347;
assign n_4349 =  x_1658 & ~n_4252;
assign n_4350 =  i_16 &  n_4252;
assign n_4351 = ~n_4349 & ~n_4350;
assign n_4352 =  x_1658 & ~n_4351;
assign n_4353 = ~x_1658 &  n_4351;
assign n_4354 = ~n_4352 & ~n_4353;
assign n_4355 =  x_1657 & ~n_4252;
assign n_4356 =  i_15 &  n_4252;
assign n_4357 = ~n_4355 & ~n_4356;
assign n_4358 =  x_1657 & ~n_4357;
assign n_4359 = ~x_1657 &  n_4357;
assign n_4360 = ~n_4358 & ~n_4359;
assign n_4361 =  x_1656 & ~n_4252;
assign n_4362 =  i_14 &  n_4252;
assign n_4363 = ~n_4361 & ~n_4362;
assign n_4364 =  x_1656 & ~n_4363;
assign n_4365 = ~x_1656 &  n_4363;
assign n_4366 = ~n_4364 & ~n_4365;
assign n_4367 =  x_1655 & ~n_4252;
assign n_4368 =  i_13 &  n_4252;
assign n_4369 = ~n_4367 & ~n_4368;
assign n_4370 =  x_1655 & ~n_4369;
assign n_4371 = ~x_1655 &  n_4369;
assign n_4372 = ~n_4370 & ~n_4371;
assign n_4373 =  x_1654 & ~n_4252;
assign n_4374 =  i_12 &  n_4252;
assign n_4375 = ~n_4373 & ~n_4374;
assign n_4376 =  x_1654 & ~n_4375;
assign n_4377 = ~x_1654 &  n_4375;
assign n_4378 = ~n_4376 & ~n_4377;
assign n_4379 =  x_1653 & ~n_4252;
assign n_4380 =  i_11 &  n_4252;
assign n_4381 = ~n_4379 & ~n_4380;
assign n_4382 =  x_1653 & ~n_4381;
assign n_4383 = ~x_1653 &  n_4381;
assign n_4384 = ~n_4382 & ~n_4383;
assign n_4385 =  x_1652 & ~n_4252;
assign n_4386 =  i_10 &  n_4252;
assign n_4387 = ~n_4385 & ~n_4386;
assign n_4388 =  x_1652 & ~n_4387;
assign n_4389 = ~x_1652 &  n_4387;
assign n_4390 = ~n_4388 & ~n_4389;
assign n_4391 =  x_1651 & ~n_4252;
assign n_4392 =  i_9 &  n_4252;
assign n_4393 = ~n_4391 & ~n_4392;
assign n_4394 =  x_1651 & ~n_4393;
assign n_4395 = ~x_1651 &  n_4393;
assign n_4396 = ~n_4394 & ~n_4395;
assign n_4397 =  x_1650 & ~n_4252;
assign n_4398 =  i_8 &  n_4252;
assign n_4399 = ~n_4397 & ~n_4398;
assign n_4400 =  x_1650 & ~n_4399;
assign n_4401 = ~x_1650 &  n_4399;
assign n_4402 = ~n_4400 & ~n_4401;
assign n_4403 =  x_1649 & ~n_4252;
assign n_4404 =  i_7 &  n_4252;
assign n_4405 = ~n_4403 & ~n_4404;
assign n_4406 =  x_1649 & ~n_4405;
assign n_4407 = ~x_1649 &  n_4405;
assign n_4408 = ~n_4406 & ~n_4407;
assign n_4409 =  x_1648 & ~n_4252;
assign n_4410 =  i_6 &  n_4252;
assign n_4411 = ~n_4409 & ~n_4410;
assign n_4412 =  x_1648 & ~n_4411;
assign n_4413 = ~x_1648 &  n_4411;
assign n_4414 = ~n_4412 & ~n_4413;
assign n_4415 =  x_1647 & ~n_4252;
assign n_4416 =  i_5 &  n_4252;
assign n_4417 = ~n_4415 & ~n_4416;
assign n_4418 =  x_1647 & ~n_4417;
assign n_4419 = ~x_1647 &  n_4417;
assign n_4420 = ~n_4418 & ~n_4419;
assign n_4421 =  x_1646 & ~n_4252;
assign n_4422 =  i_4 &  n_4252;
assign n_4423 = ~n_4421 & ~n_4422;
assign n_4424 =  x_1646 & ~n_4423;
assign n_4425 = ~x_1646 &  n_4423;
assign n_4426 = ~n_4424 & ~n_4425;
assign n_4427 =  x_1645 & ~n_4252;
assign n_4428 =  i_3 &  n_4252;
assign n_4429 = ~n_4427 & ~n_4428;
assign n_4430 =  x_1645 & ~n_4429;
assign n_4431 = ~x_1645 &  n_4429;
assign n_4432 = ~n_4430 & ~n_4431;
assign n_4433 =  x_1644 & ~n_4252;
assign n_4434 =  i_2 &  n_4252;
assign n_4435 = ~n_4433 & ~n_4434;
assign n_4436 =  x_1644 & ~n_4435;
assign n_4437 = ~x_1644 &  n_4435;
assign n_4438 = ~n_4436 & ~n_4437;
assign n_4439 =  x_1643 & ~n_4252;
assign n_4440 =  i_1 &  n_4252;
assign n_4441 = ~n_4439 & ~n_4440;
assign n_4442 =  x_1643 & ~n_4441;
assign n_4443 = ~x_1643 &  n_4441;
assign n_4444 = ~n_4442 & ~n_4443;
assign n_4445 =  n_389 &  n_1178;
assign n_4446 =  n_3 &  n_4445;
assign n_4447 =  x_1642 & ~n_4446;
assign n_4448 =  x_106 &  n_4446;
assign n_4449 = ~n_4447 & ~n_4448;
assign n_4450 =  x_1642 & ~n_4449;
assign n_4451 = ~x_1642 &  n_4449;
assign n_4452 = ~n_4450 & ~n_4451;
assign n_4453 =  x_1641 & ~n_4446;
assign n_4454 =  x_105 &  n_4446;
assign n_4455 = ~n_4453 & ~n_4454;
assign n_4456 =  x_1641 & ~n_4455;
assign n_4457 = ~x_1641 &  n_4455;
assign n_4458 = ~n_4456 & ~n_4457;
assign n_4459 =  x_1640 & ~n_4446;
assign n_4460 =  x_104 &  n_4446;
assign n_4461 = ~n_4459 & ~n_4460;
assign n_4462 =  x_1640 & ~n_4461;
assign n_4463 = ~x_1640 &  n_4461;
assign n_4464 = ~n_4462 & ~n_4463;
assign n_4465 =  x_1639 & ~n_4446;
assign n_4466 =  x_103 &  n_4446;
assign n_4467 = ~n_4465 & ~n_4466;
assign n_4468 =  x_1639 & ~n_4467;
assign n_4469 = ~x_1639 &  n_4467;
assign n_4470 = ~n_4468 & ~n_4469;
assign n_4471 =  x_1638 & ~n_4446;
assign n_4472 =  x_102 &  n_4446;
assign n_4473 = ~n_4471 & ~n_4472;
assign n_4474 =  x_1638 & ~n_4473;
assign n_4475 = ~x_1638 &  n_4473;
assign n_4476 = ~n_4474 & ~n_4475;
assign n_4477 =  x_1637 & ~n_4446;
assign n_4478 =  x_101 &  n_4446;
assign n_4479 = ~n_4477 & ~n_4478;
assign n_4480 =  x_1637 & ~n_4479;
assign n_4481 = ~x_1637 &  n_4479;
assign n_4482 = ~n_4480 & ~n_4481;
assign n_4483 =  x_1636 & ~n_4446;
assign n_4484 =  x_100 &  n_4446;
assign n_4485 = ~n_4483 & ~n_4484;
assign n_4486 =  x_1636 & ~n_4485;
assign n_4487 = ~x_1636 &  n_4485;
assign n_4488 = ~n_4486 & ~n_4487;
assign n_4489 =  x_1635 & ~n_4446;
assign n_4490 =  x_99 &  n_4446;
assign n_4491 = ~n_4489 & ~n_4490;
assign n_4492 =  x_1635 & ~n_4491;
assign n_4493 = ~x_1635 &  n_4491;
assign n_4494 = ~n_4492 & ~n_4493;
assign n_4495 =  x_1634 & ~n_4446;
assign n_4496 =  x_98 &  n_4446;
assign n_4497 = ~n_4495 & ~n_4496;
assign n_4498 =  x_1634 & ~n_4497;
assign n_4499 = ~x_1634 &  n_4497;
assign n_4500 = ~n_4498 & ~n_4499;
assign n_4501 =  x_1633 & ~n_4446;
assign n_4502 =  x_97 &  n_4446;
assign n_4503 = ~n_4501 & ~n_4502;
assign n_4504 =  x_1633 & ~n_4503;
assign n_4505 = ~x_1633 &  n_4503;
assign n_4506 = ~n_4504 & ~n_4505;
assign n_4507 =  x_1632 & ~n_4446;
assign n_4508 =  x_96 &  n_4446;
assign n_4509 = ~n_4507 & ~n_4508;
assign n_4510 =  x_1632 & ~n_4509;
assign n_4511 = ~x_1632 &  n_4509;
assign n_4512 = ~n_4510 & ~n_4511;
assign n_4513 =  x_1631 & ~n_4446;
assign n_4514 =  x_95 &  n_4446;
assign n_4515 = ~n_4513 & ~n_4514;
assign n_4516 =  x_1631 & ~n_4515;
assign n_4517 = ~x_1631 &  n_4515;
assign n_4518 = ~n_4516 & ~n_4517;
assign n_4519 =  x_1630 & ~n_4446;
assign n_4520 =  x_94 &  n_4446;
assign n_4521 = ~n_4519 & ~n_4520;
assign n_4522 =  x_1630 & ~n_4521;
assign n_4523 = ~x_1630 &  n_4521;
assign n_4524 = ~n_4522 & ~n_4523;
assign n_4525 =  x_1629 & ~n_4446;
assign n_4526 =  x_93 &  n_4446;
assign n_4527 = ~n_4525 & ~n_4526;
assign n_4528 =  x_1629 & ~n_4527;
assign n_4529 = ~x_1629 &  n_4527;
assign n_4530 = ~n_4528 & ~n_4529;
assign n_4531 =  x_1628 & ~n_4446;
assign n_4532 =  x_92 &  n_4446;
assign n_4533 = ~n_4531 & ~n_4532;
assign n_4534 =  x_1628 & ~n_4533;
assign n_4535 = ~x_1628 &  n_4533;
assign n_4536 = ~n_4534 & ~n_4535;
assign n_4537 =  x_1627 & ~n_4446;
assign n_4538 =  x_91 &  n_4446;
assign n_4539 = ~n_4537 & ~n_4538;
assign n_4540 =  x_1627 & ~n_4539;
assign n_4541 = ~x_1627 &  n_4539;
assign n_4542 = ~n_4540 & ~n_4541;
assign n_4543 =  x_1626 & ~n_4446;
assign n_4544 =  x_90 &  n_4446;
assign n_4545 = ~n_4543 & ~n_4544;
assign n_4546 =  x_1626 & ~n_4545;
assign n_4547 = ~x_1626 &  n_4545;
assign n_4548 = ~n_4546 & ~n_4547;
assign n_4549 =  x_1625 & ~n_4446;
assign n_4550 =  x_89 &  n_4446;
assign n_4551 = ~n_4549 & ~n_4550;
assign n_4552 =  x_1625 & ~n_4551;
assign n_4553 = ~x_1625 &  n_4551;
assign n_4554 = ~n_4552 & ~n_4553;
assign n_4555 =  x_1624 & ~n_4446;
assign n_4556 =  x_88 &  n_4446;
assign n_4557 = ~n_4555 & ~n_4556;
assign n_4558 =  x_1624 & ~n_4557;
assign n_4559 = ~x_1624 &  n_4557;
assign n_4560 = ~n_4558 & ~n_4559;
assign n_4561 =  x_1623 & ~n_4446;
assign n_4562 =  x_87 &  n_4446;
assign n_4563 = ~n_4561 & ~n_4562;
assign n_4564 =  x_1623 & ~n_4563;
assign n_4565 = ~x_1623 &  n_4563;
assign n_4566 = ~n_4564 & ~n_4565;
assign n_4567 =  x_1622 & ~n_4446;
assign n_4568 =  x_86 &  n_4446;
assign n_4569 = ~n_4567 & ~n_4568;
assign n_4570 =  x_1622 & ~n_4569;
assign n_4571 = ~x_1622 &  n_4569;
assign n_4572 = ~n_4570 & ~n_4571;
assign n_4573 =  x_1621 & ~n_4446;
assign n_4574 =  x_85 &  n_4446;
assign n_4575 = ~n_4573 & ~n_4574;
assign n_4576 =  x_1621 & ~n_4575;
assign n_4577 = ~x_1621 &  n_4575;
assign n_4578 = ~n_4576 & ~n_4577;
assign n_4579 =  x_1620 & ~n_4446;
assign n_4580 =  x_84 &  n_4446;
assign n_4581 = ~n_4579 & ~n_4580;
assign n_4582 =  x_1620 & ~n_4581;
assign n_4583 = ~x_1620 &  n_4581;
assign n_4584 = ~n_4582 & ~n_4583;
assign n_4585 =  x_1619 & ~n_4446;
assign n_4586 =  x_83 &  n_4446;
assign n_4587 = ~n_4585 & ~n_4586;
assign n_4588 =  x_1619 & ~n_4587;
assign n_4589 = ~x_1619 &  n_4587;
assign n_4590 = ~n_4588 & ~n_4589;
assign n_4591 =  x_1618 & ~n_4446;
assign n_4592 =  x_82 &  n_4446;
assign n_4593 = ~n_4591 & ~n_4592;
assign n_4594 =  x_1618 & ~n_4593;
assign n_4595 = ~x_1618 &  n_4593;
assign n_4596 = ~n_4594 & ~n_4595;
assign n_4597 =  x_1617 & ~n_4446;
assign n_4598 =  x_81 &  n_4446;
assign n_4599 = ~n_4597 & ~n_4598;
assign n_4600 =  x_1617 & ~n_4599;
assign n_4601 = ~x_1617 &  n_4599;
assign n_4602 = ~n_4600 & ~n_4601;
assign n_4603 =  x_1616 & ~n_4446;
assign n_4604 =  x_80 &  n_4446;
assign n_4605 = ~n_4603 & ~n_4604;
assign n_4606 =  x_1616 & ~n_4605;
assign n_4607 = ~x_1616 &  n_4605;
assign n_4608 = ~n_4606 & ~n_4607;
assign n_4609 =  x_1615 & ~n_4446;
assign n_4610 =  x_79 &  n_4446;
assign n_4611 = ~n_4609 & ~n_4610;
assign n_4612 =  x_1615 & ~n_4611;
assign n_4613 = ~x_1615 &  n_4611;
assign n_4614 = ~n_4612 & ~n_4613;
assign n_4615 =  x_1614 & ~n_4446;
assign n_4616 =  x_78 &  n_4446;
assign n_4617 = ~n_4615 & ~n_4616;
assign n_4618 =  x_1614 & ~n_4617;
assign n_4619 = ~x_1614 &  n_4617;
assign n_4620 = ~n_4618 & ~n_4619;
assign n_4621 =  x_1613 & ~n_4446;
assign n_4622 =  x_77 &  n_4446;
assign n_4623 = ~n_4621 & ~n_4622;
assign n_4624 =  x_1613 & ~n_4623;
assign n_4625 = ~x_1613 &  n_4623;
assign n_4626 = ~n_4624 & ~n_4625;
assign n_4627 =  x_1612 & ~n_4446;
assign n_4628 =  x_76 &  n_4446;
assign n_4629 = ~n_4627 & ~n_4628;
assign n_4630 =  x_1612 & ~n_4629;
assign n_4631 = ~x_1612 &  n_4629;
assign n_4632 = ~n_4630 & ~n_4631;
assign n_4633 =  x_1611 & ~n_4446;
assign n_4634 =  x_75 &  n_4446;
assign n_4635 = ~n_4633 & ~n_4634;
assign n_4636 =  x_1611 & ~n_4635;
assign n_4637 = ~x_1611 &  n_4635;
assign n_4638 = ~n_4636 & ~n_4637;
assign n_4639 =  n_186 &  n_1179;
assign n_4640 =  x_1610 & ~n_4639;
assign n_4641 =  i_32 &  n_4639;
assign n_4642 = ~n_4640 & ~n_4641;
assign n_4643 =  x_1610 & ~n_4642;
assign n_4644 = ~x_1610 &  n_4642;
assign n_4645 = ~n_4643 & ~n_4644;
assign n_4646 =  x_1609 & ~n_4639;
assign n_4647 =  i_31 &  n_4639;
assign n_4648 = ~n_4646 & ~n_4647;
assign n_4649 =  x_1609 & ~n_4648;
assign n_4650 = ~x_1609 &  n_4648;
assign n_4651 = ~n_4649 & ~n_4650;
assign n_4652 =  x_1608 & ~n_4639;
assign n_4653 =  i_30 &  n_4639;
assign n_4654 = ~n_4652 & ~n_4653;
assign n_4655 =  x_1608 & ~n_4654;
assign n_4656 = ~x_1608 &  n_4654;
assign n_4657 = ~n_4655 & ~n_4656;
assign n_4658 =  x_1607 & ~n_4639;
assign n_4659 =  i_29 &  n_4639;
assign n_4660 = ~n_4658 & ~n_4659;
assign n_4661 =  x_1607 & ~n_4660;
assign n_4662 = ~x_1607 &  n_4660;
assign n_4663 = ~n_4661 & ~n_4662;
assign n_4664 =  x_1606 & ~n_4639;
assign n_4665 =  i_28 &  n_4639;
assign n_4666 = ~n_4664 & ~n_4665;
assign n_4667 =  x_1606 & ~n_4666;
assign n_4668 = ~x_1606 &  n_4666;
assign n_4669 = ~n_4667 & ~n_4668;
assign n_4670 =  x_1605 & ~n_4639;
assign n_4671 =  i_27 &  n_4639;
assign n_4672 = ~n_4670 & ~n_4671;
assign n_4673 =  x_1605 & ~n_4672;
assign n_4674 = ~x_1605 &  n_4672;
assign n_4675 = ~n_4673 & ~n_4674;
assign n_4676 =  x_1604 & ~n_4639;
assign n_4677 =  i_26 &  n_4639;
assign n_4678 = ~n_4676 & ~n_4677;
assign n_4679 =  x_1604 & ~n_4678;
assign n_4680 = ~x_1604 &  n_4678;
assign n_4681 = ~n_4679 & ~n_4680;
assign n_4682 =  x_1603 & ~n_4639;
assign n_4683 =  i_25 &  n_4639;
assign n_4684 = ~n_4682 & ~n_4683;
assign n_4685 =  x_1603 & ~n_4684;
assign n_4686 = ~x_1603 &  n_4684;
assign n_4687 = ~n_4685 & ~n_4686;
assign n_4688 =  x_1602 & ~n_4639;
assign n_4689 =  i_24 &  n_4639;
assign n_4690 = ~n_4688 & ~n_4689;
assign n_4691 =  x_1602 & ~n_4690;
assign n_4692 = ~x_1602 &  n_4690;
assign n_4693 = ~n_4691 & ~n_4692;
assign n_4694 =  x_1601 & ~n_4639;
assign n_4695 =  i_23 &  n_4639;
assign n_4696 = ~n_4694 & ~n_4695;
assign n_4697 =  x_1601 & ~n_4696;
assign n_4698 = ~x_1601 &  n_4696;
assign n_4699 = ~n_4697 & ~n_4698;
assign n_4700 =  x_1600 & ~n_4639;
assign n_4701 =  i_22 &  n_4639;
assign n_4702 = ~n_4700 & ~n_4701;
assign n_4703 =  x_1600 & ~n_4702;
assign n_4704 = ~x_1600 &  n_4702;
assign n_4705 = ~n_4703 & ~n_4704;
assign n_4706 =  x_1599 & ~n_4639;
assign n_4707 =  i_21 &  n_4639;
assign n_4708 = ~n_4706 & ~n_4707;
assign n_4709 =  x_1599 & ~n_4708;
assign n_4710 = ~x_1599 &  n_4708;
assign n_4711 = ~n_4709 & ~n_4710;
assign n_4712 =  x_1598 & ~n_4639;
assign n_4713 =  i_20 &  n_4639;
assign n_4714 = ~n_4712 & ~n_4713;
assign n_4715 =  x_1598 & ~n_4714;
assign n_4716 = ~x_1598 &  n_4714;
assign n_4717 = ~n_4715 & ~n_4716;
assign n_4718 =  x_1597 & ~n_4639;
assign n_4719 =  i_19 &  n_4639;
assign n_4720 = ~n_4718 & ~n_4719;
assign n_4721 =  x_1597 & ~n_4720;
assign n_4722 = ~x_1597 &  n_4720;
assign n_4723 = ~n_4721 & ~n_4722;
assign n_4724 =  x_1596 & ~n_4639;
assign n_4725 =  i_18 &  n_4639;
assign n_4726 = ~n_4724 & ~n_4725;
assign n_4727 =  x_1596 & ~n_4726;
assign n_4728 = ~x_1596 &  n_4726;
assign n_4729 = ~n_4727 & ~n_4728;
assign n_4730 =  x_1595 & ~n_4639;
assign n_4731 =  i_17 &  n_4639;
assign n_4732 = ~n_4730 & ~n_4731;
assign n_4733 =  x_1595 & ~n_4732;
assign n_4734 = ~x_1595 &  n_4732;
assign n_4735 = ~n_4733 & ~n_4734;
assign n_4736 =  x_1594 & ~n_4639;
assign n_4737 =  i_16 &  n_4639;
assign n_4738 = ~n_4736 & ~n_4737;
assign n_4739 =  x_1594 & ~n_4738;
assign n_4740 = ~x_1594 &  n_4738;
assign n_4741 = ~n_4739 & ~n_4740;
assign n_4742 =  x_1593 & ~n_4639;
assign n_4743 =  i_15 &  n_4639;
assign n_4744 = ~n_4742 & ~n_4743;
assign n_4745 =  x_1593 & ~n_4744;
assign n_4746 = ~x_1593 &  n_4744;
assign n_4747 = ~n_4745 & ~n_4746;
assign n_4748 =  x_1592 & ~n_4639;
assign n_4749 =  i_14 &  n_4639;
assign n_4750 = ~n_4748 & ~n_4749;
assign n_4751 =  x_1592 & ~n_4750;
assign n_4752 = ~x_1592 &  n_4750;
assign n_4753 = ~n_4751 & ~n_4752;
assign n_4754 =  x_1591 & ~n_4639;
assign n_4755 =  i_13 &  n_4639;
assign n_4756 = ~n_4754 & ~n_4755;
assign n_4757 =  x_1591 & ~n_4756;
assign n_4758 = ~x_1591 &  n_4756;
assign n_4759 = ~n_4757 & ~n_4758;
assign n_4760 =  x_1590 & ~n_4639;
assign n_4761 =  i_12 &  n_4639;
assign n_4762 = ~n_4760 & ~n_4761;
assign n_4763 =  x_1590 & ~n_4762;
assign n_4764 = ~x_1590 &  n_4762;
assign n_4765 = ~n_4763 & ~n_4764;
assign n_4766 =  x_1589 & ~n_4639;
assign n_4767 =  i_11 &  n_4639;
assign n_4768 = ~n_4766 & ~n_4767;
assign n_4769 =  x_1589 & ~n_4768;
assign n_4770 = ~x_1589 &  n_4768;
assign n_4771 = ~n_4769 & ~n_4770;
assign n_4772 =  x_1588 & ~n_4639;
assign n_4773 =  i_10 &  n_4639;
assign n_4774 = ~n_4772 & ~n_4773;
assign n_4775 =  x_1588 & ~n_4774;
assign n_4776 = ~x_1588 &  n_4774;
assign n_4777 = ~n_4775 & ~n_4776;
assign n_4778 =  x_1587 & ~n_4639;
assign n_4779 =  i_9 &  n_4639;
assign n_4780 = ~n_4778 & ~n_4779;
assign n_4781 =  x_1587 & ~n_4780;
assign n_4782 = ~x_1587 &  n_4780;
assign n_4783 = ~n_4781 & ~n_4782;
assign n_4784 =  x_1586 & ~n_4639;
assign n_4785 =  i_8 &  n_4639;
assign n_4786 = ~n_4784 & ~n_4785;
assign n_4787 =  x_1586 & ~n_4786;
assign n_4788 = ~x_1586 &  n_4786;
assign n_4789 = ~n_4787 & ~n_4788;
assign n_4790 =  x_1585 & ~n_4639;
assign n_4791 =  i_7 &  n_4639;
assign n_4792 = ~n_4790 & ~n_4791;
assign n_4793 =  x_1585 & ~n_4792;
assign n_4794 = ~x_1585 &  n_4792;
assign n_4795 = ~n_4793 & ~n_4794;
assign n_4796 =  x_1584 & ~n_4639;
assign n_4797 =  i_6 &  n_4639;
assign n_4798 = ~n_4796 & ~n_4797;
assign n_4799 =  x_1584 & ~n_4798;
assign n_4800 = ~x_1584 &  n_4798;
assign n_4801 = ~n_4799 & ~n_4800;
assign n_4802 =  x_1583 & ~n_4639;
assign n_4803 =  i_5 &  n_4639;
assign n_4804 = ~n_4802 & ~n_4803;
assign n_4805 =  x_1583 & ~n_4804;
assign n_4806 = ~x_1583 &  n_4804;
assign n_4807 = ~n_4805 & ~n_4806;
assign n_4808 =  x_1582 & ~n_4639;
assign n_4809 =  i_4 &  n_4639;
assign n_4810 = ~n_4808 & ~n_4809;
assign n_4811 =  x_1582 & ~n_4810;
assign n_4812 = ~x_1582 &  n_4810;
assign n_4813 = ~n_4811 & ~n_4812;
assign n_4814 =  x_1581 & ~n_4639;
assign n_4815 =  i_3 &  n_4639;
assign n_4816 = ~n_4814 & ~n_4815;
assign n_4817 =  x_1581 & ~n_4816;
assign n_4818 = ~x_1581 &  n_4816;
assign n_4819 = ~n_4817 & ~n_4818;
assign n_4820 =  x_1580 & ~n_4639;
assign n_4821 =  i_2 &  n_4639;
assign n_4822 = ~n_4820 & ~n_4821;
assign n_4823 =  x_1580 & ~n_4822;
assign n_4824 = ~x_1580 &  n_4822;
assign n_4825 = ~n_4823 & ~n_4824;
assign n_4826 =  x_1579 & ~n_4639;
assign n_4827 =  i_1 &  n_4639;
assign n_4828 = ~n_4826 & ~n_4827;
assign n_4829 =  x_1579 & ~n_4828;
assign n_4830 = ~x_1579 &  n_4828;
assign n_4831 = ~n_4829 & ~n_4830;
assign n_4832 =  x_1578 & ~n_984;
assign n_4833 = ~n_985 & ~n_4832;
assign n_4834 =  x_1578 & ~n_4833;
assign n_4835 = ~x_1578 &  n_4833;
assign n_4836 = ~n_4834 & ~n_4835;
assign n_4837 =  x_1577 & ~n_984;
assign n_4838 = ~n_991 & ~n_4837;
assign n_4839 =  x_1577 & ~n_4838;
assign n_4840 = ~x_1577 &  n_4838;
assign n_4841 = ~n_4839 & ~n_4840;
assign n_4842 =  x_1576 & ~n_984;
assign n_4843 = ~n_997 & ~n_4842;
assign n_4844 =  x_1576 & ~n_4843;
assign n_4845 = ~x_1576 &  n_4843;
assign n_4846 = ~n_4844 & ~n_4845;
assign n_4847 =  x_1575 & ~n_984;
assign n_4848 = ~n_1003 & ~n_4847;
assign n_4849 =  x_1575 & ~n_4848;
assign n_4850 = ~x_1575 &  n_4848;
assign n_4851 = ~n_4849 & ~n_4850;
assign n_4852 =  x_1574 & ~n_984;
assign n_4853 = ~n_1009 & ~n_4852;
assign n_4854 =  x_1574 & ~n_4853;
assign n_4855 = ~x_1574 &  n_4853;
assign n_4856 = ~n_4854 & ~n_4855;
assign n_4857 =  x_1573 & ~n_984;
assign n_4858 = ~n_1015 & ~n_4857;
assign n_4859 =  x_1573 & ~n_4858;
assign n_4860 = ~x_1573 &  n_4858;
assign n_4861 = ~n_4859 & ~n_4860;
assign n_4862 =  x_1572 & ~n_984;
assign n_4863 = ~n_1021 & ~n_4862;
assign n_4864 =  x_1572 & ~n_4863;
assign n_4865 = ~x_1572 &  n_4863;
assign n_4866 = ~n_4864 & ~n_4865;
assign n_4867 =  x_1571 & ~n_984;
assign n_4868 = ~n_1027 & ~n_4867;
assign n_4869 =  x_1571 & ~n_4868;
assign n_4870 = ~x_1571 &  n_4868;
assign n_4871 = ~n_4869 & ~n_4870;
assign n_4872 =  x_1570 & ~n_984;
assign n_4873 = ~n_1033 & ~n_4872;
assign n_4874 =  x_1570 & ~n_4873;
assign n_4875 = ~x_1570 &  n_4873;
assign n_4876 = ~n_4874 & ~n_4875;
assign n_4877 =  x_1569 & ~n_984;
assign n_4878 = ~n_1039 & ~n_4877;
assign n_4879 =  x_1569 & ~n_4878;
assign n_4880 = ~x_1569 &  n_4878;
assign n_4881 = ~n_4879 & ~n_4880;
assign n_4882 =  x_1568 & ~n_984;
assign n_4883 = ~n_1045 & ~n_4882;
assign n_4884 =  x_1568 & ~n_4883;
assign n_4885 = ~x_1568 &  n_4883;
assign n_4886 = ~n_4884 & ~n_4885;
assign n_4887 =  x_1567 & ~n_984;
assign n_4888 = ~n_1051 & ~n_4887;
assign n_4889 =  x_1567 & ~n_4888;
assign n_4890 = ~x_1567 &  n_4888;
assign n_4891 = ~n_4889 & ~n_4890;
assign n_4892 =  x_1566 & ~n_984;
assign n_4893 = ~n_1057 & ~n_4892;
assign n_4894 =  x_1566 & ~n_4893;
assign n_4895 = ~x_1566 &  n_4893;
assign n_4896 = ~n_4894 & ~n_4895;
assign n_4897 =  x_1565 & ~n_984;
assign n_4898 = ~n_1063 & ~n_4897;
assign n_4899 =  x_1565 & ~n_4898;
assign n_4900 = ~x_1565 &  n_4898;
assign n_4901 = ~n_4899 & ~n_4900;
assign n_4902 =  x_1564 & ~n_984;
assign n_4903 = ~n_1069 & ~n_4902;
assign n_4904 =  x_1564 & ~n_4903;
assign n_4905 = ~x_1564 &  n_4903;
assign n_4906 = ~n_4904 & ~n_4905;
assign n_4907 =  x_1563 & ~n_984;
assign n_4908 = ~n_1075 & ~n_4907;
assign n_4909 =  x_1563 & ~n_4908;
assign n_4910 = ~x_1563 &  n_4908;
assign n_4911 = ~n_4909 & ~n_4910;
assign n_4912 =  x_1562 & ~n_984;
assign n_4913 = ~n_1081 & ~n_4912;
assign n_4914 =  x_1562 & ~n_4913;
assign n_4915 = ~x_1562 &  n_4913;
assign n_4916 = ~n_4914 & ~n_4915;
assign n_4917 =  x_1561 & ~n_984;
assign n_4918 = ~n_1087 & ~n_4917;
assign n_4919 =  x_1561 & ~n_4918;
assign n_4920 = ~x_1561 &  n_4918;
assign n_4921 = ~n_4919 & ~n_4920;
assign n_4922 =  x_1560 & ~n_984;
assign n_4923 = ~n_1093 & ~n_4922;
assign n_4924 =  x_1560 & ~n_4923;
assign n_4925 = ~x_1560 &  n_4923;
assign n_4926 = ~n_4924 & ~n_4925;
assign n_4927 =  x_1559 & ~n_984;
assign n_4928 = ~n_1099 & ~n_4927;
assign n_4929 =  x_1559 & ~n_4928;
assign n_4930 = ~x_1559 &  n_4928;
assign n_4931 = ~n_4929 & ~n_4930;
assign n_4932 =  x_1558 & ~n_984;
assign n_4933 = ~n_1105 & ~n_4932;
assign n_4934 =  x_1558 & ~n_4933;
assign n_4935 = ~x_1558 &  n_4933;
assign n_4936 = ~n_4934 & ~n_4935;
assign n_4937 =  x_1557 & ~n_984;
assign n_4938 = ~n_1111 & ~n_4937;
assign n_4939 =  x_1557 & ~n_4938;
assign n_4940 = ~x_1557 &  n_4938;
assign n_4941 = ~n_4939 & ~n_4940;
assign n_4942 =  x_1556 & ~n_984;
assign n_4943 = ~n_1117 & ~n_4942;
assign n_4944 =  x_1556 & ~n_4943;
assign n_4945 = ~x_1556 &  n_4943;
assign n_4946 = ~n_4944 & ~n_4945;
assign n_4947 =  x_1555 & ~n_984;
assign n_4948 = ~n_1123 & ~n_4947;
assign n_4949 =  x_1555 & ~n_4948;
assign n_4950 = ~x_1555 &  n_4948;
assign n_4951 = ~n_4949 & ~n_4950;
assign n_4952 =  x_1554 & ~n_984;
assign n_4953 = ~n_1129 & ~n_4952;
assign n_4954 =  x_1554 & ~n_4953;
assign n_4955 = ~x_1554 &  n_4953;
assign n_4956 = ~n_4954 & ~n_4955;
assign n_4957 =  x_1553 & ~n_984;
assign n_4958 = ~n_1135 & ~n_4957;
assign n_4959 =  x_1553 & ~n_4958;
assign n_4960 = ~x_1553 &  n_4958;
assign n_4961 = ~n_4959 & ~n_4960;
assign n_4962 =  x_1552 & ~n_984;
assign n_4963 = ~n_1141 & ~n_4962;
assign n_4964 =  x_1552 & ~n_4963;
assign n_4965 = ~x_1552 &  n_4963;
assign n_4966 = ~n_4964 & ~n_4965;
assign n_4967 =  x_1551 & ~n_984;
assign n_4968 = ~n_1147 & ~n_4967;
assign n_4969 =  x_1551 & ~n_4968;
assign n_4970 = ~x_1551 &  n_4968;
assign n_4971 = ~n_4969 & ~n_4970;
assign n_4972 =  x_1550 & ~n_984;
assign n_4973 = ~n_1153 & ~n_4972;
assign n_4974 =  x_1550 & ~n_4973;
assign n_4975 = ~x_1550 &  n_4973;
assign n_4976 = ~n_4974 & ~n_4975;
assign n_4977 =  x_1549 & ~n_984;
assign n_4978 = ~n_1159 & ~n_4977;
assign n_4979 =  x_1549 & ~n_4978;
assign n_4980 = ~x_1549 &  n_4978;
assign n_4981 = ~n_4979 & ~n_4980;
assign n_4982 =  x_1548 & ~n_984;
assign n_4983 = ~n_1165 & ~n_4982;
assign n_4984 =  x_1548 & ~n_4983;
assign n_4985 = ~x_1548 &  n_4983;
assign n_4986 = ~n_4984 & ~n_4985;
assign n_4987 =  x_1547 & ~n_984;
assign n_4988 = ~n_1171 & ~n_4987;
assign n_4989 =  x_1547 & ~n_4988;
assign n_4990 = ~x_1547 &  n_4988;
assign n_4991 = ~n_4989 & ~n_4990;
assign n_4992 =  x_41 &  x_42;
assign n_4993 =  n_184 &  n_4992;
assign n_4994 =  n_4993 &  n_1179;
assign n_4995 =  x_1546 & ~n_4994;
assign n_4996 =  i_32 &  n_4994;
assign n_4997 = ~n_4995 & ~n_4996;
assign n_4998 =  x_1546 & ~n_4997;
assign n_4999 = ~x_1546 &  n_4997;
assign n_5000 = ~n_4998 & ~n_4999;
assign n_5001 =  x_1545 & ~n_4994;
assign n_5002 =  i_31 &  n_4994;
assign n_5003 = ~n_5001 & ~n_5002;
assign n_5004 =  x_1545 & ~n_5003;
assign n_5005 = ~x_1545 &  n_5003;
assign n_5006 = ~n_5004 & ~n_5005;
assign n_5007 =  x_1544 & ~n_4994;
assign n_5008 =  i_30 &  n_4994;
assign n_5009 = ~n_5007 & ~n_5008;
assign n_5010 =  x_1544 & ~n_5009;
assign n_5011 = ~x_1544 &  n_5009;
assign n_5012 = ~n_5010 & ~n_5011;
assign n_5013 =  x_1543 & ~n_4994;
assign n_5014 =  i_29 &  n_4994;
assign n_5015 = ~n_5013 & ~n_5014;
assign n_5016 =  x_1543 & ~n_5015;
assign n_5017 = ~x_1543 &  n_5015;
assign n_5018 = ~n_5016 & ~n_5017;
assign n_5019 =  x_1542 & ~n_4994;
assign n_5020 =  i_28 &  n_4994;
assign n_5021 = ~n_5019 & ~n_5020;
assign n_5022 =  x_1542 & ~n_5021;
assign n_5023 = ~x_1542 &  n_5021;
assign n_5024 = ~n_5022 & ~n_5023;
assign n_5025 =  x_1541 & ~n_4994;
assign n_5026 =  i_27 &  n_4994;
assign n_5027 = ~n_5025 & ~n_5026;
assign n_5028 =  x_1541 & ~n_5027;
assign n_5029 = ~x_1541 &  n_5027;
assign n_5030 = ~n_5028 & ~n_5029;
assign n_5031 =  x_1540 & ~n_4994;
assign n_5032 =  i_26 &  n_4994;
assign n_5033 = ~n_5031 & ~n_5032;
assign n_5034 =  x_1540 & ~n_5033;
assign n_5035 = ~x_1540 &  n_5033;
assign n_5036 = ~n_5034 & ~n_5035;
assign n_5037 =  x_1539 & ~n_4994;
assign n_5038 =  i_25 &  n_4994;
assign n_5039 = ~n_5037 & ~n_5038;
assign n_5040 =  x_1539 & ~n_5039;
assign n_5041 = ~x_1539 &  n_5039;
assign n_5042 = ~n_5040 & ~n_5041;
assign n_5043 =  x_1538 & ~n_4994;
assign n_5044 =  i_24 &  n_4994;
assign n_5045 = ~n_5043 & ~n_5044;
assign n_5046 =  x_1538 & ~n_5045;
assign n_5047 = ~x_1538 &  n_5045;
assign n_5048 = ~n_5046 & ~n_5047;
assign n_5049 =  x_1537 & ~n_4994;
assign n_5050 =  i_23 &  n_4994;
assign n_5051 = ~n_5049 & ~n_5050;
assign n_5052 =  x_1537 & ~n_5051;
assign n_5053 = ~x_1537 &  n_5051;
assign n_5054 = ~n_5052 & ~n_5053;
assign n_5055 =  x_1536 & ~n_4994;
assign n_5056 =  i_22 &  n_4994;
assign n_5057 = ~n_5055 & ~n_5056;
assign n_5058 =  x_1536 & ~n_5057;
assign n_5059 = ~x_1536 &  n_5057;
assign n_5060 = ~n_5058 & ~n_5059;
assign n_5061 =  x_1535 & ~n_4994;
assign n_5062 =  i_21 &  n_4994;
assign n_5063 = ~n_5061 & ~n_5062;
assign n_5064 =  x_1535 & ~n_5063;
assign n_5065 = ~x_1535 &  n_5063;
assign n_5066 = ~n_5064 & ~n_5065;
assign n_5067 =  x_1534 & ~n_4994;
assign n_5068 =  i_20 &  n_4994;
assign n_5069 = ~n_5067 & ~n_5068;
assign n_5070 =  x_1534 & ~n_5069;
assign n_5071 = ~x_1534 &  n_5069;
assign n_5072 = ~n_5070 & ~n_5071;
assign n_5073 =  x_1533 & ~n_4994;
assign n_5074 =  i_19 &  n_4994;
assign n_5075 = ~n_5073 & ~n_5074;
assign n_5076 =  x_1533 & ~n_5075;
assign n_5077 = ~x_1533 &  n_5075;
assign n_5078 = ~n_5076 & ~n_5077;
assign n_5079 =  x_1532 & ~n_4994;
assign n_5080 =  i_18 &  n_4994;
assign n_5081 = ~n_5079 & ~n_5080;
assign n_5082 =  x_1532 & ~n_5081;
assign n_5083 = ~x_1532 &  n_5081;
assign n_5084 = ~n_5082 & ~n_5083;
assign n_5085 =  x_1531 & ~n_4994;
assign n_5086 =  i_17 &  n_4994;
assign n_5087 = ~n_5085 & ~n_5086;
assign n_5088 =  x_1531 & ~n_5087;
assign n_5089 = ~x_1531 &  n_5087;
assign n_5090 = ~n_5088 & ~n_5089;
assign n_5091 =  x_1530 & ~n_4994;
assign n_5092 =  i_16 &  n_4994;
assign n_5093 = ~n_5091 & ~n_5092;
assign n_5094 =  x_1530 & ~n_5093;
assign n_5095 = ~x_1530 &  n_5093;
assign n_5096 = ~n_5094 & ~n_5095;
assign n_5097 =  x_1529 & ~n_4994;
assign n_5098 =  i_15 &  n_4994;
assign n_5099 = ~n_5097 & ~n_5098;
assign n_5100 =  x_1529 & ~n_5099;
assign n_5101 = ~x_1529 &  n_5099;
assign n_5102 = ~n_5100 & ~n_5101;
assign n_5103 =  x_1528 & ~n_4994;
assign n_5104 =  i_14 &  n_4994;
assign n_5105 = ~n_5103 & ~n_5104;
assign n_5106 =  x_1528 & ~n_5105;
assign n_5107 = ~x_1528 &  n_5105;
assign n_5108 = ~n_5106 & ~n_5107;
assign n_5109 =  x_1527 & ~n_4994;
assign n_5110 =  i_13 &  n_4994;
assign n_5111 = ~n_5109 & ~n_5110;
assign n_5112 =  x_1527 & ~n_5111;
assign n_5113 = ~x_1527 &  n_5111;
assign n_5114 = ~n_5112 & ~n_5113;
assign n_5115 =  x_1526 & ~n_4994;
assign n_5116 =  i_12 &  n_4994;
assign n_5117 = ~n_5115 & ~n_5116;
assign n_5118 =  x_1526 & ~n_5117;
assign n_5119 = ~x_1526 &  n_5117;
assign n_5120 = ~n_5118 & ~n_5119;
assign n_5121 =  x_1525 & ~n_4994;
assign n_5122 =  i_11 &  n_4994;
assign n_5123 = ~n_5121 & ~n_5122;
assign n_5124 =  x_1525 & ~n_5123;
assign n_5125 = ~x_1525 &  n_5123;
assign n_5126 = ~n_5124 & ~n_5125;
assign n_5127 =  x_1524 & ~n_4994;
assign n_5128 =  i_10 &  n_4994;
assign n_5129 = ~n_5127 & ~n_5128;
assign n_5130 =  x_1524 & ~n_5129;
assign n_5131 = ~x_1524 &  n_5129;
assign n_5132 = ~n_5130 & ~n_5131;
assign n_5133 =  x_1523 & ~n_4994;
assign n_5134 =  i_9 &  n_4994;
assign n_5135 = ~n_5133 & ~n_5134;
assign n_5136 =  x_1523 & ~n_5135;
assign n_5137 = ~x_1523 &  n_5135;
assign n_5138 = ~n_5136 & ~n_5137;
assign n_5139 =  x_1522 & ~n_4994;
assign n_5140 =  i_8 &  n_4994;
assign n_5141 = ~n_5139 & ~n_5140;
assign n_5142 =  x_1522 & ~n_5141;
assign n_5143 = ~x_1522 &  n_5141;
assign n_5144 = ~n_5142 & ~n_5143;
assign n_5145 =  x_1521 & ~n_4994;
assign n_5146 =  i_7 &  n_4994;
assign n_5147 = ~n_5145 & ~n_5146;
assign n_5148 =  x_1521 & ~n_5147;
assign n_5149 = ~x_1521 &  n_5147;
assign n_5150 = ~n_5148 & ~n_5149;
assign n_5151 =  x_1520 & ~n_4994;
assign n_5152 =  i_6 &  n_4994;
assign n_5153 = ~n_5151 & ~n_5152;
assign n_5154 =  x_1520 & ~n_5153;
assign n_5155 = ~x_1520 &  n_5153;
assign n_5156 = ~n_5154 & ~n_5155;
assign n_5157 =  x_1519 & ~n_4994;
assign n_5158 =  i_5 &  n_4994;
assign n_5159 = ~n_5157 & ~n_5158;
assign n_5160 =  x_1519 & ~n_5159;
assign n_5161 = ~x_1519 &  n_5159;
assign n_5162 = ~n_5160 & ~n_5161;
assign n_5163 =  x_1518 & ~n_4994;
assign n_5164 =  i_4 &  n_4994;
assign n_5165 = ~n_5163 & ~n_5164;
assign n_5166 =  x_1518 & ~n_5165;
assign n_5167 = ~x_1518 &  n_5165;
assign n_5168 = ~n_5166 & ~n_5167;
assign n_5169 =  x_1517 & ~n_4994;
assign n_5170 =  i_3 &  n_4994;
assign n_5171 = ~n_5169 & ~n_5170;
assign n_5172 =  x_1517 & ~n_5171;
assign n_5173 = ~x_1517 &  n_5171;
assign n_5174 = ~n_5172 & ~n_5173;
assign n_5175 =  x_1516 & ~n_4994;
assign n_5176 =  i_2 &  n_4994;
assign n_5177 = ~n_5175 & ~n_5176;
assign n_5178 =  x_1516 & ~n_5177;
assign n_5179 = ~x_1516 &  n_5177;
assign n_5180 = ~n_5178 & ~n_5179;
assign n_5181 =  x_1515 & ~n_4994;
assign n_5182 =  i_1 &  n_4994;
assign n_5183 = ~n_5181 & ~n_5182;
assign n_5184 =  x_1515 & ~n_5183;
assign n_5185 = ~x_1515 &  n_5183;
assign n_5186 = ~n_5184 & ~n_5185;
assign n_5187 =  x_39 &  n_3081;
assign n_5188 = ~n_1709 & ~n_5187;
assign n_5189 =  n_2 & ~n_5188;
assign n_5190 =  x_1514 & ~n_5189;
assign n_5191 =  n_1708 &  n_2302;
assign n_5192 =  n_2 &  n_5191;
assign n_5193 =  x_618 &  x_2090;
assign n_5194 = ~x_618 & ~x_2090;
assign n_5195 = ~n_5193 & ~n_5194;
assign n_5196 =  n_5192 &  n_5195;
assign n_5197 =  n_3 &  n_1709;
assign n_5198 =  x_170 &  x_2826;
assign n_5199 = ~x_170 & ~x_2826;
assign n_5200 = ~n_5198 & ~n_5199;
assign n_5201 =  n_5197 &  n_5200;
assign n_5202 = ~n_5196 & ~n_5201;
assign n_5203 = ~n_5190 &  n_5202;
assign n_5204 =  x_1514 & ~n_5203;
assign n_5205 = ~x_1514 &  n_5203;
assign n_5206 = ~n_5204 & ~n_5205;
assign n_5207 =  x_1513 & ~n_5189;
assign n_5208 = ~x_2089 & ~x_2090;
assign n_5209 =  x_2089 &  x_2090;
assign n_5210 = ~n_5208 & ~n_5209;
assign n_5211 =  x_617 &  n_5210;
assign n_5212 = ~x_617 & ~n_5210;
assign n_5213 = ~n_5211 & ~n_5212;
assign n_5214 =  n_5193 &  n_5213;
assign n_5215 = ~n_5193 & ~n_5213;
assign n_5216 =  n_5192 & ~n_5215;
assign n_5217 = ~n_5214 &  n_5216;
assign n_5218 = ~x_169 & ~x_170;
assign n_5219 =  x_169 &  x_170;
assign n_5220 = ~n_5218 & ~n_5219;
assign n_5221 =  x_2825 &  n_5220;
assign n_5222 = ~x_2825 & ~n_5220;
assign n_5223 = ~n_5221 & ~n_5222;
assign n_5224 = ~n_5198 & ~n_5223;
assign n_5225 =  n_5198 &  n_5223;
assign n_5226 =  n_5197 & ~n_5225;
assign n_5227 = ~n_5224 &  n_5226;
assign n_5228 = ~n_5217 & ~n_5227;
assign n_5229 = ~n_5207 &  n_5228;
assign n_5230 =  x_1513 & ~n_5229;
assign n_5231 = ~x_1513 &  n_5229;
assign n_5232 = ~n_5230 & ~n_5231;
assign n_5233 = ~x_2088 &  n_5208;
assign n_5234 =  x_2088 & ~n_5208;
assign n_5235 = ~n_5233 & ~n_5234;
assign n_5236 = ~x_617 &  x_2089;
assign n_5237 =  n_5193 & ~n_5236;
assign n_5238 = ~n_5237 & ~n_5211;
assign n_5239 =  n_5235 & ~n_5238;
assign n_5240 = ~n_5235 &  n_5238;
assign n_5241 = ~n_5239 & ~n_5240;
assign n_5242 = ~x_616 & ~n_5241;
assign n_5243 =  x_616 & ~n_5240;
assign n_5244 = ~n_5239 &  n_5243;
assign n_5245 =  n_5192 & ~n_5244;
assign n_5246 = ~n_5242 &  n_5245;
assign n_5247 =  x_1512 & ~n_5189;
assign n_5248 = ~x_168 &  n_5218;
assign n_5249 =  x_168 & ~n_5218;
assign n_5250 = ~n_5248 & ~n_5249;
assign n_5251 =  x_169 & ~x_2825;
assign n_5252 =  n_5198 & ~n_5251;
assign n_5253 = ~n_5252 & ~n_5221;
assign n_5254 =  n_5250 & ~n_5253;
assign n_5255 = ~n_5250 &  n_5253;
assign n_5256 = ~n_5254 & ~n_5255;
assign n_5257 = ~x_2824 & ~n_5256;
assign n_5258 =  x_2824 & ~n_5255;
assign n_5259 = ~n_5254 &  n_5258;
assign n_5260 =  n_5197 & ~n_5259;
assign n_5261 = ~n_5257 &  n_5260;
assign n_5262 = ~n_5247 & ~n_5261;
assign n_5263 = ~n_5246 &  n_5262;
assign n_5264 =  x_1512 & ~n_5263;
assign n_5265 = ~x_1512 &  n_5263;
assign n_5266 = ~n_5264 & ~n_5265;
assign n_5267 = ~x_167 &  n_5248;
assign n_5268 =  x_167 & ~n_5248;
assign n_5269 = ~n_5267 & ~n_5268;
assign n_5270 = ~n_5254 & ~n_5258;
assign n_5271 =  n_5269 & ~n_5270;
assign n_5272 = ~n_5269 &  n_5270;
assign n_5273 = ~n_5271 & ~n_5272;
assign n_5274 = ~x_2823 & ~n_5273;
assign n_5275 =  x_2823 & ~n_5272;
assign n_5276 = ~n_5271 &  n_5275;
assign n_5277 =  n_5197 & ~n_5276;
assign n_5278 = ~n_5274 &  n_5277;
assign n_5279 =  x_1511 & ~n_5189;
assign n_5280 = ~x_2087 &  n_5233;
assign n_5281 =  x_2087 & ~n_5233;
assign n_5282 = ~n_5280 & ~n_5281;
assign n_5283 = ~n_5239 & ~n_5243;
assign n_5284 =  n_5282 & ~n_5283;
assign n_5285 = ~n_5282 &  n_5283;
assign n_5286 = ~n_5284 & ~n_5285;
assign n_5287 = ~x_615 & ~n_5286;
assign n_5288 =  x_615 & ~n_5285;
assign n_5289 = ~n_5284 &  n_5288;
assign n_5290 =  n_5192 & ~n_5289;
assign n_5291 = ~n_5287 &  n_5290;
assign n_5292 = ~n_5279 & ~n_5291;
assign n_5293 = ~n_5278 &  n_5292;
assign n_5294 =  x_1511 & ~n_5293;
assign n_5295 = ~x_1511 &  n_5293;
assign n_5296 = ~n_5294 & ~n_5295;
assign n_5297 = ~x_166 &  n_5267;
assign n_5298 =  x_166 & ~n_5267;
assign n_5299 = ~n_5297 & ~n_5298;
assign n_5300 = ~n_5271 & ~n_5275;
assign n_5301 =  n_5299 & ~n_5300;
assign n_5302 = ~n_5299 &  n_5300;
assign n_5303 = ~n_5301 & ~n_5302;
assign n_5304 = ~x_2822 & ~n_5303;
assign n_5305 =  x_2822 & ~n_5302;
assign n_5306 = ~n_5301 &  n_5305;
assign n_5307 =  n_5197 & ~n_5306;
assign n_5308 = ~n_5304 &  n_5307;
assign n_5309 =  x_1510 & ~n_5189;
assign n_5310 = ~x_2086 &  n_5280;
assign n_5311 =  x_2086 & ~n_5280;
assign n_5312 = ~n_5310 & ~n_5311;
assign n_5313 = ~n_5284 & ~n_5288;
assign n_5314 =  n_5312 & ~n_5313;
assign n_5315 = ~n_5312 &  n_5313;
assign n_5316 = ~n_5314 & ~n_5315;
assign n_5317 = ~x_614 & ~n_5316;
assign n_5318 =  x_614 & ~n_5315;
assign n_5319 = ~n_5314 &  n_5318;
assign n_5320 =  n_5192 & ~n_5319;
assign n_5321 = ~n_5317 &  n_5320;
assign n_5322 = ~n_5309 & ~n_5321;
assign n_5323 = ~n_5308 &  n_5322;
assign n_5324 =  x_1510 & ~n_5323;
assign n_5325 = ~x_1510 &  n_5323;
assign n_5326 = ~n_5324 & ~n_5325;
assign n_5327 = ~x_165 &  n_5297;
assign n_5328 =  x_165 & ~n_5297;
assign n_5329 = ~n_5327 & ~n_5328;
assign n_5330 = ~n_5301 & ~n_5305;
assign n_5331 =  n_5329 & ~n_5330;
assign n_5332 = ~n_5329 &  n_5330;
assign n_5333 = ~n_5331 & ~n_5332;
assign n_5334 = ~x_2821 & ~n_5333;
assign n_5335 =  x_2821 & ~n_5332;
assign n_5336 = ~n_5331 &  n_5335;
assign n_5337 =  n_5197 & ~n_5336;
assign n_5338 = ~n_5334 &  n_5337;
assign n_5339 =  x_1509 & ~n_5189;
assign n_5340 = ~x_2085 &  n_5310;
assign n_5341 =  x_2085 & ~n_5310;
assign n_5342 = ~n_5340 & ~n_5341;
assign n_5343 = ~n_5314 & ~n_5318;
assign n_5344 =  n_5342 & ~n_5343;
assign n_5345 = ~n_5342 &  n_5343;
assign n_5346 = ~n_5344 & ~n_5345;
assign n_5347 = ~x_613 & ~n_5346;
assign n_5348 =  x_613 & ~n_5345;
assign n_5349 = ~n_5344 &  n_5348;
assign n_5350 =  n_5192 & ~n_5349;
assign n_5351 = ~n_5347 &  n_5350;
assign n_5352 = ~n_5339 & ~n_5351;
assign n_5353 = ~n_5338 &  n_5352;
assign n_5354 =  x_1509 & ~n_5353;
assign n_5355 = ~x_1509 &  n_5353;
assign n_5356 = ~n_5354 & ~n_5355;
assign n_5357 = ~x_164 &  n_5327;
assign n_5358 =  x_164 & ~n_5327;
assign n_5359 = ~n_5357 & ~n_5358;
assign n_5360 = ~n_5331 & ~n_5335;
assign n_5361 =  n_5359 & ~n_5360;
assign n_5362 = ~n_5359 &  n_5360;
assign n_5363 = ~n_5361 & ~n_5362;
assign n_5364 = ~x_2820 & ~n_5363;
assign n_5365 =  x_2820 & ~n_5362;
assign n_5366 = ~n_5361 &  n_5365;
assign n_5367 =  n_5197 & ~n_5366;
assign n_5368 = ~n_5364 &  n_5367;
assign n_5369 =  x_1508 & ~n_5189;
assign n_5370 = ~x_2084 &  n_5340;
assign n_5371 =  x_2084 & ~n_5340;
assign n_5372 = ~n_5370 & ~n_5371;
assign n_5373 = ~n_5344 & ~n_5348;
assign n_5374 =  n_5372 & ~n_5373;
assign n_5375 = ~n_5372 &  n_5373;
assign n_5376 = ~n_5374 & ~n_5375;
assign n_5377 = ~x_612 & ~n_5376;
assign n_5378 =  x_612 & ~n_5375;
assign n_5379 = ~n_5374 &  n_5378;
assign n_5380 =  n_5192 & ~n_5379;
assign n_5381 = ~n_5377 &  n_5380;
assign n_5382 = ~n_5369 & ~n_5381;
assign n_5383 = ~n_5368 &  n_5382;
assign n_5384 =  x_1508 & ~n_5383;
assign n_5385 = ~x_1508 &  n_5383;
assign n_5386 = ~n_5384 & ~n_5385;
assign n_5387 = ~x_163 &  n_5357;
assign n_5388 =  x_163 & ~n_5357;
assign n_5389 = ~n_5387 & ~n_5388;
assign n_5390 = ~n_5361 & ~n_5365;
assign n_5391 =  n_5389 & ~n_5390;
assign n_5392 = ~n_5389 &  n_5390;
assign n_5393 = ~n_5391 & ~n_5392;
assign n_5394 = ~x_2819 & ~n_5393;
assign n_5395 =  x_2819 & ~n_5392;
assign n_5396 = ~n_5391 &  n_5395;
assign n_5397 =  n_5197 & ~n_5396;
assign n_5398 = ~n_5394 &  n_5397;
assign n_5399 =  x_1507 & ~n_5189;
assign n_5400 = ~x_2083 &  n_5370;
assign n_5401 =  x_2083 & ~n_5370;
assign n_5402 = ~n_5400 & ~n_5401;
assign n_5403 = ~n_5374 & ~n_5378;
assign n_5404 =  n_5402 & ~n_5403;
assign n_5405 = ~n_5402 &  n_5403;
assign n_5406 = ~n_5404 & ~n_5405;
assign n_5407 = ~x_611 & ~n_5406;
assign n_5408 =  x_611 & ~n_5405;
assign n_5409 = ~n_5404 &  n_5408;
assign n_5410 =  n_5192 & ~n_5409;
assign n_5411 = ~n_5407 &  n_5410;
assign n_5412 = ~n_5399 & ~n_5411;
assign n_5413 = ~n_5398 &  n_5412;
assign n_5414 =  x_1507 & ~n_5413;
assign n_5415 = ~x_1507 &  n_5413;
assign n_5416 = ~n_5414 & ~n_5415;
assign n_5417 = ~x_162 &  n_5387;
assign n_5418 =  x_162 & ~n_5387;
assign n_5419 = ~n_5417 & ~n_5418;
assign n_5420 = ~n_5391 & ~n_5395;
assign n_5421 =  n_5419 & ~n_5420;
assign n_5422 = ~n_5419 &  n_5420;
assign n_5423 = ~n_5421 & ~n_5422;
assign n_5424 = ~x_2818 & ~n_5423;
assign n_5425 =  x_2818 & ~n_5422;
assign n_5426 = ~n_5421 &  n_5425;
assign n_5427 =  n_5197 & ~n_5426;
assign n_5428 = ~n_5424 &  n_5427;
assign n_5429 =  x_1506 & ~n_5189;
assign n_5430 = ~x_2082 &  n_5400;
assign n_5431 =  x_2082 & ~n_5400;
assign n_5432 = ~n_5430 & ~n_5431;
assign n_5433 = ~n_5404 & ~n_5408;
assign n_5434 =  n_5432 & ~n_5433;
assign n_5435 = ~n_5432 &  n_5433;
assign n_5436 = ~n_5434 & ~n_5435;
assign n_5437 = ~x_610 & ~n_5436;
assign n_5438 =  x_610 & ~n_5435;
assign n_5439 = ~n_5434 &  n_5438;
assign n_5440 =  n_5192 & ~n_5439;
assign n_5441 = ~n_5437 &  n_5440;
assign n_5442 = ~n_5429 & ~n_5441;
assign n_5443 = ~n_5428 &  n_5442;
assign n_5444 =  x_1506 & ~n_5443;
assign n_5445 = ~x_1506 &  n_5443;
assign n_5446 = ~n_5444 & ~n_5445;
assign n_5447 = ~x_161 &  n_5417;
assign n_5448 =  x_161 & ~n_5417;
assign n_5449 = ~n_5447 & ~n_5448;
assign n_5450 = ~n_5421 & ~n_5425;
assign n_5451 =  n_5449 & ~n_5450;
assign n_5452 = ~n_5449 &  n_5450;
assign n_5453 = ~n_5451 & ~n_5452;
assign n_5454 = ~x_2817 & ~n_5453;
assign n_5455 =  x_2817 & ~n_5452;
assign n_5456 = ~n_5451 &  n_5455;
assign n_5457 =  n_5197 & ~n_5456;
assign n_5458 = ~n_5454 &  n_5457;
assign n_5459 =  x_1505 & ~n_5189;
assign n_5460 = ~x_2081 &  n_5430;
assign n_5461 =  x_2081 & ~n_5430;
assign n_5462 = ~n_5460 & ~n_5461;
assign n_5463 = ~n_5434 & ~n_5438;
assign n_5464 =  n_5462 & ~n_5463;
assign n_5465 = ~n_5462 &  n_5463;
assign n_5466 = ~n_5464 & ~n_5465;
assign n_5467 = ~x_609 & ~n_5466;
assign n_5468 =  x_609 & ~n_5465;
assign n_5469 = ~n_5464 &  n_5468;
assign n_5470 =  n_5192 & ~n_5469;
assign n_5471 = ~n_5467 &  n_5470;
assign n_5472 = ~n_5459 & ~n_5471;
assign n_5473 = ~n_5458 &  n_5472;
assign n_5474 =  x_1505 & ~n_5473;
assign n_5475 = ~x_1505 &  n_5473;
assign n_5476 = ~n_5474 & ~n_5475;
assign n_5477 = ~x_160 &  n_5447;
assign n_5478 =  x_160 & ~n_5447;
assign n_5479 = ~n_5477 & ~n_5478;
assign n_5480 = ~n_5451 & ~n_5455;
assign n_5481 =  n_5479 & ~n_5480;
assign n_5482 = ~n_5479 &  n_5480;
assign n_5483 = ~n_5481 & ~n_5482;
assign n_5484 = ~x_2816 & ~n_5483;
assign n_5485 =  x_2816 & ~n_5482;
assign n_5486 = ~n_5481 &  n_5485;
assign n_5487 =  n_5197 & ~n_5486;
assign n_5488 = ~n_5484 &  n_5487;
assign n_5489 =  x_1504 & ~n_5189;
assign n_5490 = ~x_2080 &  n_5460;
assign n_5491 =  x_2080 & ~n_5460;
assign n_5492 = ~n_5490 & ~n_5491;
assign n_5493 = ~n_5464 & ~n_5468;
assign n_5494 =  n_5492 & ~n_5493;
assign n_5495 = ~n_5492 &  n_5493;
assign n_5496 = ~n_5494 & ~n_5495;
assign n_5497 = ~x_608 & ~n_5496;
assign n_5498 =  x_608 & ~n_5495;
assign n_5499 = ~n_5494 &  n_5498;
assign n_5500 =  n_5192 & ~n_5499;
assign n_5501 = ~n_5497 &  n_5500;
assign n_5502 = ~n_5489 & ~n_5501;
assign n_5503 = ~n_5488 &  n_5502;
assign n_5504 =  x_1504 & ~n_5503;
assign n_5505 = ~x_1504 &  n_5503;
assign n_5506 = ~n_5504 & ~n_5505;
assign n_5507 = ~x_159 &  n_5477;
assign n_5508 =  x_159 & ~n_5477;
assign n_5509 = ~n_5507 & ~n_5508;
assign n_5510 = ~n_5481 & ~n_5485;
assign n_5511 =  n_5509 & ~n_5510;
assign n_5512 = ~n_5509 &  n_5510;
assign n_5513 = ~n_5511 & ~n_5512;
assign n_5514 = ~x_2815 & ~n_5513;
assign n_5515 =  x_2815 & ~n_5512;
assign n_5516 = ~n_5511 &  n_5515;
assign n_5517 =  n_5197 & ~n_5516;
assign n_5518 = ~n_5514 &  n_5517;
assign n_5519 =  x_1503 & ~n_5189;
assign n_5520 = ~x_2079 &  n_5490;
assign n_5521 =  x_2079 & ~n_5490;
assign n_5522 = ~n_5520 & ~n_5521;
assign n_5523 = ~n_5494 & ~n_5498;
assign n_5524 =  n_5522 & ~n_5523;
assign n_5525 = ~n_5522 &  n_5523;
assign n_5526 = ~n_5524 & ~n_5525;
assign n_5527 = ~x_607 & ~n_5526;
assign n_5528 =  x_607 & ~n_5525;
assign n_5529 = ~n_5524 &  n_5528;
assign n_5530 =  n_5192 & ~n_5529;
assign n_5531 = ~n_5527 &  n_5530;
assign n_5532 = ~n_5519 & ~n_5531;
assign n_5533 = ~n_5518 &  n_5532;
assign n_5534 =  x_1503 & ~n_5533;
assign n_5535 = ~x_1503 &  n_5533;
assign n_5536 = ~n_5534 & ~n_5535;
assign n_5537 = ~x_158 &  n_5507;
assign n_5538 =  x_158 & ~n_5507;
assign n_5539 = ~n_5537 & ~n_5538;
assign n_5540 = ~n_5511 & ~n_5515;
assign n_5541 =  n_5539 & ~n_5540;
assign n_5542 = ~n_5539 &  n_5540;
assign n_5543 = ~n_5541 & ~n_5542;
assign n_5544 = ~x_2814 & ~n_5543;
assign n_5545 =  x_2814 & ~n_5542;
assign n_5546 = ~n_5541 &  n_5545;
assign n_5547 =  n_5197 & ~n_5546;
assign n_5548 = ~n_5544 &  n_5547;
assign n_5549 =  x_1502 & ~n_5189;
assign n_5550 = ~x_2078 &  n_5520;
assign n_5551 =  x_2078 & ~n_5520;
assign n_5552 = ~n_5550 & ~n_5551;
assign n_5553 = ~n_5524 & ~n_5528;
assign n_5554 =  n_5552 & ~n_5553;
assign n_5555 = ~n_5552 &  n_5553;
assign n_5556 = ~n_5554 & ~n_5555;
assign n_5557 = ~x_606 & ~n_5556;
assign n_5558 =  x_606 & ~n_5555;
assign n_5559 = ~n_5554 &  n_5558;
assign n_5560 =  n_5192 & ~n_5559;
assign n_5561 = ~n_5557 &  n_5560;
assign n_5562 = ~n_5549 & ~n_5561;
assign n_5563 = ~n_5548 &  n_5562;
assign n_5564 =  x_1502 & ~n_5563;
assign n_5565 = ~x_1502 &  n_5563;
assign n_5566 = ~n_5564 & ~n_5565;
assign n_5567 = ~x_157 &  n_5537;
assign n_5568 =  x_157 & ~n_5537;
assign n_5569 = ~n_5567 & ~n_5568;
assign n_5570 = ~n_5541 & ~n_5545;
assign n_5571 =  n_5569 & ~n_5570;
assign n_5572 = ~n_5569 &  n_5570;
assign n_5573 = ~n_5571 & ~n_5572;
assign n_5574 = ~x_2813 & ~n_5573;
assign n_5575 =  x_2813 & ~n_5572;
assign n_5576 = ~n_5571 &  n_5575;
assign n_5577 =  n_5197 & ~n_5576;
assign n_5578 = ~n_5574 &  n_5577;
assign n_5579 =  x_1501 & ~n_5189;
assign n_5580 = ~x_2077 &  n_5550;
assign n_5581 =  x_2077 & ~n_5550;
assign n_5582 = ~n_5580 & ~n_5581;
assign n_5583 = ~n_5554 & ~n_5558;
assign n_5584 =  n_5582 & ~n_5583;
assign n_5585 = ~n_5582 &  n_5583;
assign n_5586 = ~n_5584 & ~n_5585;
assign n_5587 = ~x_605 & ~n_5586;
assign n_5588 =  x_605 & ~n_5585;
assign n_5589 = ~n_5584 &  n_5588;
assign n_5590 =  n_5192 & ~n_5589;
assign n_5591 = ~n_5587 &  n_5590;
assign n_5592 = ~n_5579 & ~n_5591;
assign n_5593 = ~n_5578 &  n_5592;
assign n_5594 =  x_1501 & ~n_5593;
assign n_5595 = ~x_1501 &  n_5593;
assign n_5596 = ~n_5594 & ~n_5595;
assign n_5597 = ~x_156 &  n_5567;
assign n_5598 =  x_156 & ~n_5567;
assign n_5599 = ~n_5597 & ~n_5598;
assign n_5600 = ~n_5571 & ~n_5575;
assign n_5601 =  n_5599 & ~n_5600;
assign n_5602 = ~n_5599 &  n_5600;
assign n_5603 = ~n_5601 & ~n_5602;
assign n_5604 = ~x_2812 & ~n_5603;
assign n_5605 =  x_2812 & ~n_5602;
assign n_5606 = ~n_5601 &  n_5605;
assign n_5607 =  n_5197 & ~n_5606;
assign n_5608 = ~n_5604 &  n_5607;
assign n_5609 =  x_1500 & ~n_5189;
assign n_5610 = ~x_2076 &  n_5580;
assign n_5611 =  x_2076 & ~n_5580;
assign n_5612 = ~n_5610 & ~n_5611;
assign n_5613 = ~n_5584 & ~n_5588;
assign n_5614 =  n_5612 & ~n_5613;
assign n_5615 = ~n_5612 &  n_5613;
assign n_5616 = ~n_5614 & ~n_5615;
assign n_5617 = ~x_604 & ~n_5616;
assign n_5618 =  x_604 & ~n_5615;
assign n_5619 = ~n_5614 &  n_5618;
assign n_5620 =  n_5192 & ~n_5619;
assign n_5621 = ~n_5617 &  n_5620;
assign n_5622 = ~n_5609 & ~n_5621;
assign n_5623 = ~n_5608 &  n_5622;
assign n_5624 =  x_1500 & ~n_5623;
assign n_5625 = ~x_1500 &  n_5623;
assign n_5626 = ~n_5624 & ~n_5625;
assign n_5627 = ~x_155 &  n_5597;
assign n_5628 =  x_155 & ~n_5597;
assign n_5629 = ~n_5627 & ~n_5628;
assign n_5630 = ~n_5601 & ~n_5605;
assign n_5631 =  n_5629 & ~n_5630;
assign n_5632 = ~n_5629 &  n_5630;
assign n_5633 = ~n_5631 & ~n_5632;
assign n_5634 = ~x_2811 & ~n_5633;
assign n_5635 =  x_2811 & ~n_5632;
assign n_5636 = ~n_5631 &  n_5635;
assign n_5637 =  n_5197 & ~n_5636;
assign n_5638 = ~n_5634 &  n_5637;
assign n_5639 =  x_1499 & ~n_5189;
assign n_5640 = ~x_2075 &  n_5610;
assign n_5641 =  x_2075 & ~n_5610;
assign n_5642 = ~n_5640 & ~n_5641;
assign n_5643 = ~n_5614 & ~n_5618;
assign n_5644 =  n_5642 & ~n_5643;
assign n_5645 = ~n_5642 &  n_5643;
assign n_5646 = ~n_5644 & ~n_5645;
assign n_5647 = ~x_603 & ~n_5646;
assign n_5648 =  x_603 & ~n_5645;
assign n_5649 = ~n_5644 &  n_5648;
assign n_5650 =  n_5192 & ~n_5649;
assign n_5651 = ~n_5647 &  n_5650;
assign n_5652 = ~n_5639 & ~n_5651;
assign n_5653 = ~n_5638 &  n_5652;
assign n_5654 =  x_1499 & ~n_5653;
assign n_5655 = ~x_1499 &  n_5653;
assign n_5656 = ~n_5654 & ~n_5655;
assign n_5657 = ~x_154 &  n_5627;
assign n_5658 =  x_154 & ~n_5627;
assign n_5659 = ~n_5657 & ~n_5658;
assign n_5660 = ~n_5631 & ~n_5635;
assign n_5661 =  n_5659 & ~n_5660;
assign n_5662 = ~n_5659 &  n_5660;
assign n_5663 = ~n_5661 & ~n_5662;
assign n_5664 = ~x_2810 & ~n_5663;
assign n_5665 =  x_2810 & ~n_5662;
assign n_5666 = ~n_5661 &  n_5665;
assign n_5667 =  n_5197 & ~n_5666;
assign n_5668 = ~n_5664 &  n_5667;
assign n_5669 =  x_1498 & ~n_5189;
assign n_5670 = ~x_2074 &  n_5640;
assign n_5671 =  x_2074 & ~n_5640;
assign n_5672 = ~n_5670 & ~n_5671;
assign n_5673 = ~n_5644 & ~n_5648;
assign n_5674 =  n_5672 & ~n_5673;
assign n_5675 = ~n_5672 &  n_5673;
assign n_5676 = ~n_5674 & ~n_5675;
assign n_5677 = ~x_602 & ~n_5676;
assign n_5678 =  x_602 & ~n_5675;
assign n_5679 = ~n_5674 &  n_5678;
assign n_5680 =  n_5192 & ~n_5679;
assign n_5681 = ~n_5677 &  n_5680;
assign n_5682 = ~n_5669 & ~n_5681;
assign n_5683 = ~n_5668 &  n_5682;
assign n_5684 =  x_1498 & ~n_5683;
assign n_5685 = ~x_1498 &  n_5683;
assign n_5686 = ~n_5684 & ~n_5685;
assign n_5687 = ~x_153 &  n_5657;
assign n_5688 =  x_153 & ~n_5657;
assign n_5689 = ~n_5687 & ~n_5688;
assign n_5690 = ~n_5661 & ~n_5665;
assign n_5691 =  n_5689 & ~n_5690;
assign n_5692 = ~n_5689 &  n_5690;
assign n_5693 = ~n_5691 & ~n_5692;
assign n_5694 = ~x_2809 & ~n_5693;
assign n_5695 =  x_2809 & ~n_5692;
assign n_5696 = ~n_5691 &  n_5695;
assign n_5697 =  n_5197 & ~n_5696;
assign n_5698 = ~n_5694 &  n_5697;
assign n_5699 =  x_1497 & ~n_5189;
assign n_5700 = ~x_2073 &  n_5670;
assign n_5701 =  x_2073 & ~n_5670;
assign n_5702 = ~n_5700 & ~n_5701;
assign n_5703 = ~n_5674 & ~n_5678;
assign n_5704 =  n_5702 & ~n_5703;
assign n_5705 = ~n_5702 &  n_5703;
assign n_5706 = ~n_5704 & ~n_5705;
assign n_5707 = ~x_601 & ~n_5706;
assign n_5708 =  x_601 & ~n_5705;
assign n_5709 = ~n_5704 &  n_5708;
assign n_5710 =  n_5192 & ~n_5709;
assign n_5711 = ~n_5707 &  n_5710;
assign n_5712 = ~n_5699 & ~n_5711;
assign n_5713 = ~n_5698 &  n_5712;
assign n_5714 =  x_1497 & ~n_5713;
assign n_5715 = ~x_1497 &  n_5713;
assign n_5716 = ~n_5714 & ~n_5715;
assign n_5717 = ~x_152 &  n_5687;
assign n_5718 =  x_152 & ~n_5687;
assign n_5719 = ~n_5717 & ~n_5718;
assign n_5720 = ~n_5691 & ~n_5695;
assign n_5721 =  n_5719 & ~n_5720;
assign n_5722 = ~n_5719 &  n_5720;
assign n_5723 = ~n_5721 & ~n_5722;
assign n_5724 = ~x_2808 & ~n_5723;
assign n_5725 =  x_2808 & ~n_5722;
assign n_5726 = ~n_5721 &  n_5725;
assign n_5727 =  n_5197 & ~n_5726;
assign n_5728 = ~n_5724 &  n_5727;
assign n_5729 =  x_1496 & ~n_5189;
assign n_5730 = ~x_2072 &  n_5700;
assign n_5731 =  x_2072 & ~n_5700;
assign n_5732 = ~n_5730 & ~n_5731;
assign n_5733 = ~n_5704 & ~n_5708;
assign n_5734 =  n_5732 & ~n_5733;
assign n_5735 = ~n_5732 &  n_5733;
assign n_5736 = ~n_5734 & ~n_5735;
assign n_5737 = ~x_600 & ~n_5736;
assign n_5738 =  x_600 & ~n_5735;
assign n_5739 = ~n_5734 &  n_5738;
assign n_5740 =  n_5192 & ~n_5739;
assign n_5741 = ~n_5737 &  n_5740;
assign n_5742 = ~n_5729 & ~n_5741;
assign n_5743 = ~n_5728 &  n_5742;
assign n_5744 =  x_1496 & ~n_5743;
assign n_5745 = ~x_1496 &  n_5743;
assign n_5746 = ~n_5744 & ~n_5745;
assign n_5747 = ~x_151 &  n_5717;
assign n_5748 =  x_151 & ~n_5717;
assign n_5749 = ~n_5747 & ~n_5748;
assign n_5750 = ~n_5721 & ~n_5725;
assign n_5751 =  n_5749 & ~n_5750;
assign n_5752 = ~n_5749 &  n_5750;
assign n_5753 = ~n_5751 & ~n_5752;
assign n_5754 = ~x_2807 & ~n_5753;
assign n_5755 =  x_2807 & ~n_5752;
assign n_5756 = ~n_5751 &  n_5755;
assign n_5757 =  n_5197 & ~n_5756;
assign n_5758 = ~n_5754 &  n_5757;
assign n_5759 =  x_1495 & ~n_5189;
assign n_5760 = ~x_2071 &  n_5730;
assign n_5761 =  x_2071 & ~n_5730;
assign n_5762 = ~n_5760 & ~n_5761;
assign n_5763 = ~n_5734 & ~n_5738;
assign n_5764 =  n_5762 & ~n_5763;
assign n_5765 = ~n_5762 &  n_5763;
assign n_5766 = ~n_5764 & ~n_5765;
assign n_5767 = ~x_599 & ~n_5766;
assign n_5768 =  x_599 & ~n_5765;
assign n_5769 = ~n_5764 &  n_5768;
assign n_5770 =  n_5192 & ~n_5769;
assign n_5771 = ~n_5767 &  n_5770;
assign n_5772 = ~n_5759 & ~n_5771;
assign n_5773 = ~n_5758 &  n_5772;
assign n_5774 =  x_1495 & ~n_5773;
assign n_5775 = ~x_1495 &  n_5773;
assign n_5776 = ~n_5774 & ~n_5775;
assign n_5777 = ~x_150 &  n_5747;
assign n_5778 =  x_150 & ~n_5747;
assign n_5779 = ~n_5777 & ~n_5778;
assign n_5780 = ~n_5751 & ~n_5755;
assign n_5781 =  n_5779 & ~n_5780;
assign n_5782 = ~n_5779 &  n_5780;
assign n_5783 = ~n_5781 & ~n_5782;
assign n_5784 = ~x_2806 & ~n_5783;
assign n_5785 =  x_2806 & ~n_5782;
assign n_5786 = ~n_5781 &  n_5785;
assign n_5787 =  n_5197 & ~n_5786;
assign n_5788 = ~n_5784 &  n_5787;
assign n_5789 =  x_1494 & ~n_5189;
assign n_5790 = ~x_2070 &  n_5760;
assign n_5791 =  x_2070 & ~n_5760;
assign n_5792 = ~n_5790 & ~n_5791;
assign n_5793 = ~n_5764 & ~n_5768;
assign n_5794 =  n_5792 & ~n_5793;
assign n_5795 = ~n_5792 &  n_5793;
assign n_5796 = ~n_5794 & ~n_5795;
assign n_5797 = ~x_598 & ~n_5796;
assign n_5798 =  x_598 & ~n_5795;
assign n_5799 = ~n_5794 &  n_5798;
assign n_5800 =  n_5192 & ~n_5799;
assign n_5801 = ~n_5797 &  n_5800;
assign n_5802 = ~n_5789 & ~n_5801;
assign n_5803 = ~n_5788 &  n_5802;
assign n_5804 =  x_1494 & ~n_5803;
assign n_5805 = ~x_1494 &  n_5803;
assign n_5806 = ~n_5804 & ~n_5805;
assign n_5807 = ~x_149 &  n_5777;
assign n_5808 =  x_149 & ~n_5777;
assign n_5809 = ~n_5807 & ~n_5808;
assign n_5810 = ~n_5781 & ~n_5785;
assign n_5811 =  n_5809 & ~n_5810;
assign n_5812 = ~n_5809 &  n_5810;
assign n_5813 = ~n_5811 & ~n_5812;
assign n_5814 = ~x_2805 & ~n_5813;
assign n_5815 =  x_2805 & ~n_5812;
assign n_5816 = ~n_5811 &  n_5815;
assign n_5817 =  n_5197 & ~n_5816;
assign n_5818 = ~n_5814 &  n_5817;
assign n_5819 =  x_1493 & ~n_5189;
assign n_5820 = ~x_2069 &  n_5790;
assign n_5821 =  x_2069 & ~n_5790;
assign n_5822 = ~n_5820 & ~n_5821;
assign n_5823 = ~n_5794 & ~n_5798;
assign n_5824 =  n_5822 & ~n_5823;
assign n_5825 = ~n_5822 &  n_5823;
assign n_5826 = ~n_5824 & ~n_5825;
assign n_5827 = ~x_597 & ~n_5826;
assign n_5828 =  x_597 & ~n_5825;
assign n_5829 = ~n_5824 &  n_5828;
assign n_5830 =  n_5192 & ~n_5829;
assign n_5831 = ~n_5827 &  n_5830;
assign n_5832 = ~n_5819 & ~n_5831;
assign n_5833 = ~n_5818 &  n_5832;
assign n_5834 =  x_1493 & ~n_5833;
assign n_5835 = ~x_1493 &  n_5833;
assign n_5836 = ~n_5834 & ~n_5835;
assign n_5837 = ~x_148 &  n_5807;
assign n_5838 =  x_148 & ~n_5807;
assign n_5839 = ~n_5837 & ~n_5838;
assign n_5840 = ~n_5811 & ~n_5815;
assign n_5841 =  n_5839 & ~n_5840;
assign n_5842 = ~n_5839 &  n_5840;
assign n_5843 = ~n_5841 & ~n_5842;
assign n_5844 = ~x_2804 & ~n_5843;
assign n_5845 =  x_2804 & ~n_5842;
assign n_5846 = ~n_5841 &  n_5845;
assign n_5847 =  n_5197 & ~n_5846;
assign n_5848 = ~n_5844 &  n_5847;
assign n_5849 =  x_1492 & ~n_5189;
assign n_5850 = ~x_2068 &  n_5820;
assign n_5851 =  x_2068 & ~n_5820;
assign n_5852 = ~n_5850 & ~n_5851;
assign n_5853 = ~n_5824 & ~n_5828;
assign n_5854 =  n_5852 & ~n_5853;
assign n_5855 = ~n_5852 &  n_5853;
assign n_5856 = ~n_5854 & ~n_5855;
assign n_5857 = ~x_596 & ~n_5856;
assign n_5858 =  x_596 & ~n_5855;
assign n_5859 = ~n_5854 &  n_5858;
assign n_5860 =  n_5192 & ~n_5859;
assign n_5861 = ~n_5857 &  n_5860;
assign n_5862 = ~n_5849 & ~n_5861;
assign n_5863 = ~n_5848 &  n_5862;
assign n_5864 =  x_1492 & ~n_5863;
assign n_5865 = ~x_1492 &  n_5863;
assign n_5866 = ~n_5864 & ~n_5865;
assign n_5867 = ~x_147 &  n_5837;
assign n_5868 =  x_147 & ~n_5837;
assign n_5869 = ~n_5867 & ~n_5868;
assign n_5870 = ~n_5841 & ~n_5845;
assign n_5871 =  n_5869 & ~n_5870;
assign n_5872 = ~n_5869 &  n_5870;
assign n_5873 = ~n_5871 & ~n_5872;
assign n_5874 = ~x_2803 & ~n_5873;
assign n_5875 =  x_2803 & ~n_5872;
assign n_5876 = ~n_5871 &  n_5875;
assign n_5877 =  n_5197 & ~n_5876;
assign n_5878 = ~n_5874 &  n_5877;
assign n_5879 =  x_1491 & ~n_5189;
assign n_5880 = ~x_2067 &  n_5850;
assign n_5881 =  x_2067 & ~n_5850;
assign n_5882 = ~n_5880 & ~n_5881;
assign n_5883 = ~n_5854 & ~n_5858;
assign n_5884 =  n_5882 & ~n_5883;
assign n_5885 = ~n_5882 &  n_5883;
assign n_5886 = ~n_5884 & ~n_5885;
assign n_5887 = ~x_595 & ~n_5886;
assign n_5888 =  x_595 & ~n_5885;
assign n_5889 = ~n_5884 &  n_5888;
assign n_5890 =  n_5192 & ~n_5889;
assign n_5891 = ~n_5887 &  n_5890;
assign n_5892 = ~n_5879 & ~n_5891;
assign n_5893 = ~n_5878 &  n_5892;
assign n_5894 =  x_1491 & ~n_5893;
assign n_5895 = ~x_1491 &  n_5893;
assign n_5896 = ~n_5894 & ~n_5895;
assign n_5897 = ~x_146 &  n_5867;
assign n_5898 =  x_146 & ~n_5867;
assign n_5899 = ~n_5897 & ~n_5898;
assign n_5900 = ~n_5871 & ~n_5875;
assign n_5901 =  n_5899 & ~n_5900;
assign n_5902 = ~n_5899 &  n_5900;
assign n_5903 = ~n_5901 & ~n_5902;
assign n_5904 = ~x_2802 & ~n_5903;
assign n_5905 =  x_2802 & ~n_5902;
assign n_5906 = ~n_5901 &  n_5905;
assign n_5907 =  n_5197 & ~n_5906;
assign n_5908 = ~n_5904 &  n_5907;
assign n_5909 =  x_1490 & ~n_5189;
assign n_5910 = ~x_2066 &  n_5880;
assign n_5911 =  x_2066 & ~n_5880;
assign n_5912 = ~n_5910 & ~n_5911;
assign n_5913 = ~n_5884 & ~n_5888;
assign n_5914 =  n_5912 & ~n_5913;
assign n_5915 = ~n_5912 &  n_5913;
assign n_5916 = ~n_5914 & ~n_5915;
assign n_5917 = ~x_594 & ~n_5916;
assign n_5918 =  x_594 & ~n_5915;
assign n_5919 = ~n_5914 &  n_5918;
assign n_5920 =  n_5192 & ~n_5919;
assign n_5921 = ~n_5917 &  n_5920;
assign n_5922 = ~n_5909 & ~n_5921;
assign n_5923 = ~n_5908 &  n_5922;
assign n_5924 =  x_1490 & ~n_5923;
assign n_5925 = ~x_1490 &  n_5923;
assign n_5926 = ~n_5924 & ~n_5925;
assign n_5927 = ~x_145 &  n_5897;
assign n_5928 =  x_145 & ~n_5897;
assign n_5929 = ~n_5927 & ~n_5928;
assign n_5930 = ~n_5901 & ~n_5905;
assign n_5931 =  n_5929 & ~n_5930;
assign n_5932 = ~n_5929 &  n_5930;
assign n_5933 = ~n_5931 & ~n_5932;
assign n_5934 = ~x_2801 & ~n_5933;
assign n_5935 =  x_2801 & ~n_5932;
assign n_5936 = ~n_5931 &  n_5935;
assign n_5937 =  n_5197 & ~n_5936;
assign n_5938 = ~n_5934 &  n_5937;
assign n_5939 =  x_1489 & ~n_5189;
assign n_5940 = ~x_2065 &  n_5910;
assign n_5941 =  x_2065 & ~n_5910;
assign n_5942 = ~n_5940 & ~n_5941;
assign n_5943 = ~n_5914 & ~n_5918;
assign n_5944 =  n_5942 & ~n_5943;
assign n_5945 = ~n_5942 &  n_5943;
assign n_5946 = ~n_5944 & ~n_5945;
assign n_5947 = ~x_593 & ~n_5946;
assign n_5948 =  x_593 & ~n_5945;
assign n_5949 = ~n_5944 &  n_5948;
assign n_5950 =  n_5192 & ~n_5949;
assign n_5951 = ~n_5947 &  n_5950;
assign n_5952 = ~n_5939 & ~n_5951;
assign n_5953 = ~n_5938 &  n_5952;
assign n_5954 =  x_1489 & ~n_5953;
assign n_5955 = ~x_1489 &  n_5953;
assign n_5956 = ~n_5954 & ~n_5955;
assign n_5957 = ~x_144 &  n_5927;
assign n_5958 =  x_144 & ~n_5927;
assign n_5959 = ~n_5957 & ~n_5958;
assign n_5960 = ~n_5931 & ~n_5935;
assign n_5961 =  n_5959 & ~n_5960;
assign n_5962 = ~n_5959 &  n_5960;
assign n_5963 = ~n_5961 & ~n_5962;
assign n_5964 = ~x_2800 & ~n_5963;
assign n_5965 =  x_2800 & ~n_5962;
assign n_5966 = ~n_5961 &  n_5965;
assign n_5967 =  n_5197 & ~n_5966;
assign n_5968 = ~n_5964 &  n_5967;
assign n_5969 =  x_1488 & ~n_5189;
assign n_5970 = ~x_2064 &  n_5940;
assign n_5971 =  x_2064 & ~n_5940;
assign n_5972 = ~n_5970 & ~n_5971;
assign n_5973 = ~n_5944 & ~n_5948;
assign n_5974 =  n_5972 & ~n_5973;
assign n_5975 = ~n_5972 &  n_5973;
assign n_5976 = ~n_5974 & ~n_5975;
assign n_5977 = ~x_592 & ~n_5976;
assign n_5978 =  x_592 & ~n_5975;
assign n_5979 = ~n_5974 &  n_5978;
assign n_5980 =  n_5192 & ~n_5979;
assign n_5981 = ~n_5977 &  n_5980;
assign n_5982 = ~n_5969 & ~n_5981;
assign n_5983 = ~n_5968 &  n_5982;
assign n_5984 =  x_1488 & ~n_5983;
assign n_5985 = ~x_1488 &  n_5983;
assign n_5986 = ~n_5984 & ~n_5985;
assign n_5987 = ~x_143 &  n_5957;
assign n_5988 =  x_143 & ~n_5957;
assign n_5989 = ~n_5987 & ~n_5988;
assign n_5990 = ~n_5961 & ~n_5965;
assign n_5991 =  n_5989 & ~n_5990;
assign n_5992 = ~n_5989 &  n_5990;
assign n_5993 = ~n_5991 & ~n_5992;
assign n_5994 = ~x_2799 & ~n_5993;
assign n_5995 =  x_2799 & ~n_5992;
assign n_5996 = ~n_5991 &  n_5995;
assign n_5997 =  n_5197 & ~n_5996;
assign n_5998 = ~n_5994 &  n_5997;
assign n_5999 =  x_1487 & ~n_5189;
assign n_6000 = ~x_2063 &  n_5970;
assign n_6001 =  x_2063 & ~n_5970;
assign n_6002 = ~n_6000 & ~n_6001;
assign n_6003 = ~n_5974 & ~n_5978;
assign n_6004 =  n_6002 & ~n_6003;
assign n_6005 = ~n_6002 &  n_6003;
assign n_6006 = ~n_6004 & ~n_6005;
assign n_6007 = ~x_591 & ~n_6006;
assign n_6008 =  x_591 & ~n_6005;
assign n_6009 = ~n_6004 &  n_6008;
assign n_6010 =  n_5192 & ~n_6009;
assign n_6011 = ~n_6007 &  n_6010;
assign n_6012 = ~n_5999 & ~n_6011;
assign n_6013 = ~n_5998 &  n_6012;
assign n_6014 =  x_1487 & ~n_6013;
assign n_6015 = ~x_1487 &  n_6013;
assign n_6016 = ~n_6014 & ~n_6015;
assign n_6017 = ~x_142 &  n_5987;
assign n_6018 =  x_142 & ~n_5987;
assign n_6019 = ~n_6017 & ~n_6018;
assign n_6020 = ~n_5991 & ~n_5995;
assign n_6021 =  n_6019 & ~n_6020;
assign n_6022 = ~n_6019 &  n_6020;
assign n_6023 = ~n_6021 & ~n_6022;
assign n_6024 = ~x_2798 & ~n_6023;
assign n_6025 =  x_2798 & ~n_6022;
assign n_6026 = ~n_6021 &  n_6025;
assign n_6027 =  n_5197 & ~n_6026;
assign n_6028 = ~n_6024 &  n_6027;
assign n_6029 =  x_1486 & ~n_5189;
assign n_6030 = ~x_2062 &  n_6000;
assign n_6031 =  x_2062 & ~n_6000;
assign n_6032 = ~n_6030 & ~n_6031;
assign n_6033 = ~n_6004 & ~n_6008;
assign n_6034 =  n_6032 & ~n_6033;
assign n_6035 = ~n_6032 &  n_6033;
assign n_6036 = ~n_6034 & ~n_6035;
assign n_6037 = ~x_590 & ~n_6036;
assign n_6038 =  x_590 & ~n_6035;
assign n_6039 = ~n_6034 &  n_6038;
assign n_6040 =  n_5192 & ~n_6039;
assign n_6041 = ~n_6037 &  n_6040;
assign n_6042 = ~n_6029 & ~n_6041;
assign n_6043 = ~n_6028 &  n_6042;
assign n_6044 =  x_1486 & ~n_6043;
assign n_6045 = ~x_1486 &  n_6043;
assign n_6046 = ~n_6044 & ~n_6045;
assign n_6047 = ~x_141 &  n_6017;
assign n_6048 =  x_141 & ~n_6017;
assign n_6049 = ~n_6047 & ~n_6048;
assign n_6050 = ~n_6021 & ~n_6025;
assign n_6051 =  n_6049 & ~n_6050;
assign n_6052 = ~n_6049 &  n_6050;
assign n_6053 = ~n_6051 & ~n_6052;
assign n_6054 = ~x_2797 & ~n_6053;
assign n_6055 =  x_2797 & ~n_6052;
assign n_6056 = ~n_6051 &  n_6055;
assign n_6057 =  n_5197 & ~n_6056;
assign n_6058 = ~n_6054 &  n_6057;
assign n_6059 =  x_1485 & ~n_5189;
assign n_6060 = ~x_2061 &  n_6030;
assign n_6061 =  x_2061 & ~n_6030;
assign n_6062 = ~n_6060 & ~n_6061;
assign n_6063 = ~n_6034 & ~n_6038;
assign n_6064 =  n_6062 & ~n_6063;
assign n_6065 = ~n_6062 &  n_6063;
assign n_6066 = ~n_6064 & ~n_6065;
assign n_6067 = ~x_589 & ~n_6066;
assign n_6068 =  x_589 & ~n_6065;
assign n_6069 = ~n_6064 &  n_6068;
assign n_6070 =  n_5192 & ~n_6069;
assign n_6071 = ~n_6067 &  n_6070;
assign n_6072 = ~n_6059 & ~n_6071;
assign n_6073 = ~n_6058 &  n_6072;
assign n_6074 =  x_1485 & ~n_6073;
assign n_6075 = ~x_1485 &  n_6073;
assign n_6076 = ~n_6074 & ~n_6075;
assign n_6077 = ~x_140 &  n_6047;
assign n_6078 =  x_140 & ~n_6047;
assign n_6079 = ~n_6077 & ~n_6078;
assign n_6080 = ~n_6051 & ~n_6055;
assign n_6081 =  n_6079 & ~n_6080;
assign n_6082 = ~n_6079 &  n_6080;
assign n_6083 = ~n_6081 & ~n_6082;
assign n_6084 = ~x_2796 & ~n_6083;
assign n_6085 =  x_2796 & ~n_6082;
assign n_6086 = ~n_6081 &  n_6085;
assign n_6087 =  n_5197 & ~n_6086;
assign n_6088 = ~n_6084 &  n_6087;
assign n_6089 =  x_1484 & ~n_5189;
assign n_6090 = ~x_2060 &  n_6060;
assign n_6091 =  x_2060 & ~n_6060;
assign n_6092 = ~n_6090 & ~n_6091;
assign n_6093 = ~n_6064 & ~n_6068;
assign n_6094 =  n_6092 & ~n_6093;
assign n_6095 = ~n_6092 &  n_6093;
assign n_6096 = ~n_6094 & ~n_6095;
assign n_6097 = ~x_588 & ~n_6096;
assign n_6098 =  x_588 & ~n_6095;
assign n_6099 = ~n_6094 &  n_6098;
assign n_6100 =  n_5192 & ~n_6099;
assign n_6101 = ~n_6097 &  n_6100;
assign n_6102 = ~n_6089 & ~n_6101;
assign n_6103 = ~n_6088 &  n_6102;
assign n_6104 =  x_1484 & ~n_6103;
assign n_6105 = ~x_1484 &  n_6103;
assign n_6106 = ~n_6104 & ~n_6105;
assign n_6107 = ~n_6094 & ~n_6098;
assign n_6108 =  x_587 & ~x_2059;
assign n_6109 = ~x_587 &  x_2059;
assign n_6110 = ~n_6108 & ~n_6109;
assign n_6111 =  n_6090 &  n_6110;
assign n_6112 = ~n_6090 & ~n_6110;
assign n_6113 = ~n_6111 & ~n_6112;
assign n_6114 =  n_6107 & ~n_6113;
assign n_6115 = ~n_6107 &  n_6113;
assign n_6116 =  n_5192 & ~n_6115;
assign n_6117 = ~n_6114 &  n_6116;
assign n_6118 =  x_1483 & ~n_5189;
assign n_6119 = ~n_6081 & ~n_6085;
assign n_6120 =  x_139 & ~x_2795;
assign n_6121 = ~x_139 &  x_2795;
assign n_6122 = ~n_6120 & ~n_6121;
assign n_6123 =  n_6077 &  n_6122;
assign n_6124 = ~n_6077 & ~n_6122;
assign n_6125 = ~n_6123 & ~n_6124;
assign n_6126 =  n_6119 & ~n_6125;
assign n_6127 = ~n_6119 &  n_6125;
assign n_6128 =  n_5197 & ~n_6127;
assign n_6129 = ~n_6126 &  n_6128;
assign n_6130 = ~n_6118 & ~n_6129;
assign n_6131 = ~n_6117 &  n_6130;
assign n_6132 =  x_1483 & ~n_6131;
assign n_6133 = ~x_1483 &  n_6131;
assign n_6134 = ~n_6132 & ~n_6133;
assign n_6135 =  n_2100 &  n_1178;
assign n_6136 =  n_1905 &  n_6135;
assign n_6137 = ~x_42 &  n_6136;
assign n_6138 =  x_1482 & ~n_6137;
assign n_6139 =  i_32 &  n_6137;
assign n_6140 = ~n_6138 & ~n_6139;
assign n_6141 =  x_1482 & ~n_6140;
assign n_6142 = ~x_1482 &  n_6140;
assign n_6143 = ~n_6141 & ~n_6142;
assign n_6144 =  x_1481 & ~n_6137;
assign n_6145 =  i_31 &  n_6137;
assign n_6146 = ~n_6144 & ~n_6145;
assign n_6147 =  x_1481 & ~n_6146;
assign n_6148 = ~x_1481 &  n_6146;
assign n_6149 = ~n_6147 & ~n_6148;
assign n_6150 =  x_1480 & ~n_6137;
assign n_6151 =  i_30 &  n_6137;
assign n_6152 = ~n_6150 & ~n_6151;
assign n_6153 =  x_1480 & ~n_6152;
assign n_6154 = ~x_1480 &  n_6152;
assign n_6155 = ~n_6153 & ~n_6154;
assign n_6156 =  x_1479 & ~n_6137;
assign n_6157 =  i_29 &  n_6137;
assign n_6158 = ~n_6156 & ~n_6157;
assign n_6159 =  x_1479 & ~n_6158;
assign n_6160 = ~x_1479 &  n_6158;
assign n_6161 = ~n_6159 & ~n_6160;
assign n_6162 =  x_1478 & ~n_6137;
assign n_6163 =  i_28 &  n_6137;
assign n_6164 = ~n_6162 & ~n_6163;
assign n_6165 =  x_1478 & ~n_6164;
assign n_6166 = ~x_1478 &  n_6164;
assign n_6167 = ~n_6165 & ~n_6166;
assign n_6168 =  x_1477 & ~n_6137;
assign n_6169 =  i_27 &  n_6137;
assign n_6170 = ~n_6168 & ~n_6169;
assign n_6171 =  x_1477 & ~n_6170;
assign n_6172 = ~x_1477 &  n_6170;
assign n_6173 = ~n_6171 & ~n_6172;
assign n_6174 =  x_1476 & ~n_6137;
assign n_6175 =  i_26 &  n_6137;
assign n_6176 = ~n_6174 & ~n_6175;
assign n_6177 =  x_1476 & ~n_6176;
assign n_6178 = ~x_1476 &  n_6176;
assign n_6179 = ~n_6177 & ~n_6178;
assign n_6180 =  x_1475 & ~n_6137;
assign n_6181 =  i_25 &  n_6137;
assign n_6182 = ~n_6180 & ~n_6181;
assign n_6183 =  x_1475 & ~n_6182;
assign n_6184 = ~x_1475 &  n_6182;
assign n_6185 = ~n_6183 & ~n_6184;
assign n_6186 =  x_1474 & ~n_6137;
assign n_6187 =  i_24 &  n_6137;
assign n_6188 = ~n_6186 & ~n_6187;
assign n_6189 =  x_1474 & ~n_6188;
assign n_6190 = ~x_1474 &  n_6188;
assign n_6191 = ~n_6189 & ~n_6190;
assign n_6192 =  x_1473 & ~n_6137;
assign n_6193 =  i_23 &  n_6137;
assign n_6194 = ~n_6192 & ~n_6193;
assign n_6195 =  x_1473 & ~n_6194;
assign n_6196 = ~x_1473 &  n_6194;
assign n_6197 = ~n_6195 & ~n_6196;
assign n_6198 =  x_1472 & ~n_6137;
assign n_6199 =  i_22 &  n_6137;
assign n_6200 = ~n_6198 & ~n_6199;
assign n_6201 =  x_1472 & ~n_6200;
assign n_6202 = ~x_1472 &  n_6200;
assign n_6203 = ~n_6201 & ~n_6202;
assign n_6204 =  x_1471 & ~n_6137;
assign n_6205 =  i_21 &  n_6137;
assign n_6206 = ~n_6204 & ~n_6205;
assign n_6207 =  x_1471 & ~n_6206;
assign n_6208 = ~x_1471 &  n_6206;
assign n_6209 = ~n_6207 & ~n_6208;
assign n_6210 =  x_1470 & ~n_6137;
assign n_6211 =  i_20 &  n_6137;
assign n_6212 = ~n_6210 & ~n_6211;
assign n_6213 =  x_1470 & ~n_6212;
assign n_6214 = ~x_1470 &  n_6212;
assign n_6215 = ~n_6213 & ~n_6214;
assign n_6216 =  x_1469 & ~n_6137;
assign n_6217 =  i_19 &  n_6137;
assign n_6218 = ~n_6216 & ~n_6217;
assign n_6219 =  x_1469 & ~n_6218;
assign n_6220 = ~x_1469 &  n_6218;
assign n_6221 = ~n_6219 & ~n_6220;
assign n_6222 =  x_1468 & ~n_6137;
assign n_6223 =  i_18 &  n_6137;
assign n_6224 = ~n_6222 & ~n_6223;
assign n_6225 =  x_1468 & ~n_6224;
assign n_6226 = ~x_1468 &  n_6224;
assign n_6227 = ~n_6225 & ~n_6226;
assign n_6228 =  x_1467 & ~n_6137;
assign n_6229 =  i_17 &  n_6137;
assign n_6230 = ~n_6228 & ~n_6229;
assign n_6231 =  x_1467 & ~n_6230;
assign n_6232 = ~x_1467 &  n_6230;
assign n_6233 = ~n_6231 & ~n_6232;
assign n_6234 =  x_1466 & ~n_6137;
assign n_6235 =  i_16 &  n_6137;
assign n_6236 = ~n_6234 & ~n_6235;
assign n_6237 =  x_1466 & ~n_6236;
assign n_6238 = ~x_1466 &  n_6236;
assign n_6239 = ~n_6237 & ~n_6238;
assign n_6240 =  x_1465 & ~n_6137;
assign n_6241 =  i_15 &  n_6137;
assign n_6242 = ~n_6240 & ~n_6241;
assign n_6243 =  x_1465 & ~n_6242;
assign n_6244 = ~x_1465 &  n_6242;
assign n_6245 = ~n_6243 & ~n_6244;
assign n_6246 =  x_1464 & ~n_6137;
assign n_6247 =  i_14 &  n_6137;
assign n_6248 = ~n_6246 & ~n_6247;
assign n_6249 =  x_1464 & ~n_6248;
assign n_6250 = ~x_1464 &  n_6248;
assign n_6251 = ~n_6249 & ~n_6250;
assign n_6252 =  x_1463 & ~n_6137;
assign n_6253 =  i_13 &  n_6137;
assign n_6254 = ~n_6252 & ~n_6253;
assign n_6255 =  x_1463 & ~n_6254;
assign n_6256 = ~x_1463 &  n_6254;
assign n_6257 = ~n_6255 & ~n_6256;
assign n_6258 =  x_1462 & ~n_6137;
assign n_6259 =  i_12 &  n_6137;
assign n_6260 = ~n_6258 & ~n_6259;
assign n_6261 =  x_1462 & ~n_6260;
assign n_6262 = ~x_1462 &  n_6260;
assign n_6263 = ~n_6261 & ~n_6262;
assign n_6264 =  x_1461 & ~n_6137;
assign n_6265 =  i_11 &  n_6137;
assign n_6266 = ~n_6264 & ~n_6265;
assign n_6267 =  x_1461 & ~n_6266;
assign n_6268 = ~x_1461 &  n_6266;
assign n_6269 = ~n_6267 & ~n_6268;
assign n_6270 =  x_1460 & ~n_6137;
assign n_6271 =  i_10 &  n_6137;
assign n_6272 = ~n_6270 & ~n_6271;
assign n_6273 =  x_1460 & ~n_6272;
assign n_6274 = ~x_1460 &  n_6272;
assign n_6275 = ~n_6273 & ~n_6274;
assign n_6276 =  x_1459 & ~n_6137;
assign n_6277 =  i_9 &  n_6137;
assign n_6278 = ~n_6276 & ~n_6277;
assign n_6279 =  x_1459 & ~n_6278;
assign n_6280 = ~x_1459 &  n_6278;
assign n_6281 = ~n_6279 & ~n_6280;
assign n_6282 =  x_1458 & ~n_6137;
assign n_6283 =  i_8 &  n_6137;
assign n_6284 = ~n_6282 & ~n_6283;
assign n_6285 =  x_1458 & ~n_6284;
assign n_6286 = ~x_1458 &  n_6284;
assign n_6287 = ~n_6285 & ~n_6286;
assign n_6288 =  x_1457 & ~n_6137;
assign n_6289 =  i_7 &  n_6137;
assign n_6290 = ~n_6288 & ~n_6289;
assign n_6291 =  x_1457 & ~n_6290;
assign n_6292 = ~x_1457 &  n_6290;
assign n_6293 = ~n_6291 & ~n_6292;
assign n_6294 =  x_1456 & ~n_6137;
assign n_6295 =  i_6 &  n_6137;
assign n_6296 = ~n_6294 & ~n_6295;
assign n_6297 =  x_1456 & ~n_6296;
assign n_6298 = ~x_1456 &  n_6296;
assign n_6299 = ~n_6297 & ~n_6298;
assign n_6300 =  x_1455 & ~n_6137;
assign n_6301 =  i_5 &  n_6137;
assign n_6302 = ~n_6300 & ~n_6301;
assign n_6303 =  x_1455 & ~n_6302;
assign n_6304 = ~x_1455 &  n_6302;
assign n_6305 = ~n_6303 & ~n_6304;
assign n_6306 =  x_1454 & ~n_6137;
assign n_6307 =  i_4 &  n_6137;
assign n_6308 = ~n_6306 & ~n_6307;
assign n_6309 =  x_1454 & ~n_6308;
assign n_6310 = ~x_1454 &  n_6308;
assign n_6311 = ~n_6309 & ~n_6310;
assign n_6312 =  x_1453 & ~n_6137;
assign n_6313 =  i_3 &  n_6137;
assign n_6314 = ~n_6312 & ~n_6313;
assign n_6315 =  x_1453 & ~n_6314;
assign n_6316 = ~x_1453 &  n_6314;
assign n_6317 = ~n_6315 & ~n_6316;
assign n_6318 =  x_1452 & ~n_6137;
assign n_6319 =  i_2 &  n_6137;
assign n_6320 = ~n_6318 & ~n_6319;
assign n_6321 =  x_1452 & ~n_6320;
assign n_6322 = ~x_1452 &  n_6320;
assign n_6323 = ~n_6321 & ~n_6322;
assign n_6324 =  x_1451 & ~n_6137;
assign n_6325 =  i_1 &  n_6137;
assign n_6326 = ~n_6324 & ~n_6325;
assign n_6327 =  x_1451 & ~n_6326;
assign n_6328 = ~x_1451 &  n_6326;
assign n_6329 = ~n_6327 & ~n_6328;
assign n_6330 = ~x_37 &  n_1903;
assign n_6331 =  n_6330 &  n_3861;
assign n_6332 =  x_39 &  n_6135;
assign n_6333 = ~n_6331 & ~n_6332;
assign n_6334 =  n_2 & ~n_6333;
assign n_6335 =  x_1450 & ~n_6334;
assign n_6336 =  i_32 &  n_6334;
assign n_6337 = ~n_6335 & ~n_6336;
assign n_6338 =  x_1450 & ~n_6337;
assign n_6339 = ~x_1450 &  n_6337;
assign n_6340 = ~n_6338 & ~n_6339;
assign n_6341 =  x_1449 & ~n_6334;
assign n_6342 =  i_31 &  n_6334;
assign n_6343 = ~n_6341 & ~n_6342;
assign n_6344 =  x_1449 & ~n_6343;
assign n_6345 = ~x_1449 &  n_6343;
assign n_6346 = ~n_6344 & ~n_6345;
assign n_6347 =  x_1448 & ~n_6334;
assign n_6348 =  i_30 &  n_6334;
assign n_6349 = ~n_6347 & ~n_6348;
assign n_6350 =  x_1448 & ~n_6349;
assign n_6351 = ~x_1448 &  n_6349;
assign n_6352 = ~n_6350 & ~n_6351;
assign n_6353 =  x_1447 & ~n_6334;
assign n_6354 =  i_29 &  n_6334;
assign n_6355 = ~n_6353 & ~n_6354;
assign n_6356 =  x_1447 & ~n_6355;
assign n_6357 = ~x_1447 &  n_6355;
assign n_6358 = ~n_6356 & ~n_6357;
assign n_6359 =  x_1446 & ~n_6334;
assign n_6360 =  i_28 &  n_6334;
assign n_6361 = ~n_6359 & ~n_6360;
assign n_6362 =  x_1446 & ~n_6361;
assign n_6363 = ~x_1446 &  n_6361;
assign n_6364 = ~n_6362 & ~n_6363;
assign n_6365 =  x_1445 & ~n_6334;
assign n_6366 =  i_27 &  n_6334;
assign n_6367 = ~n_6365 & ~n_6366;
assign n_6368 =  x_1445 & ~n_6367;
assign n_6369 = ~x_1445 &  n_6367;
assign n_6370 = ~n_6368 & ~n_6369;
assign n_6371 =  x_1444 & ~n_6334;
assign n_6372 =  i_26 &  n_6334;
assign n_6373 = ~n_6371 & ~n_6372;
assign n_6374 =  x_1444 & ~n_6373;
assign n_6375 = ~x_1444 &  n_6373;
assign n_6376 = ~n_6374 & ~n_6375;
assign n_6377 =  x_1443 & ~n_6334;
assign n_6378 =  i_25 &  n_6334;
assign n_6379 = ~n_6377 & ~n_6378;
assign n_6380 =  x_1443 & ~n_6379;
assign n_6381 = ~x_1443 &  n_6379;
assign n_6382 = ~n_6380 & ~n_6381;
assign n_6383 =  x_1442 & ~n_6334;
assign n_6384 =  i_24 &  n_6334;
assign n_6385 = ~n_6383 & ~n_6384;
assign n_6386 =  x_1442 & ~n_6385;
assign n_6387 = ~x_1442 &  n_6385;
assign n_6388 = ~n_6386 & ~n_6387;
assign n_6389 =  x_1441 & ~n_6334;
assign n_6390 =  i_23 &  n_6334;
assign n_6391 = ~n_6389 & ~n_6390;
assign n_6392 =  x_1441 & ~n_6391;
assign n_6393 = ~x_1441 &  n_6391;
assign n_6394 = ~n_6392 & ~n_6393;
assign n_6395 =  x_1440 & ~n_6334;
assign n_6396 =  i_22 &  n_6334;
assign n_6397 = ~n_6395 & ~n_6396;
assign n_6398 =  x_1440 & ~n_6397;
assign n_6399 = ~x_1440 &  n_6397;
assign n_6400 = ~n_6398 & ~n_6399;
assign n_6401 =  x_1439 & ~n_6334;
assign n_6402 =  i_21 &  n_6334;
assign n_6403 = ~n_6401 & ~n_6402;
assign n_6404 =  x_1439 & ~n_6403;
assign n_6405 = ~x_1439 &  n_6403;
assign n_6406 = ~n_6404 & ~n_6405;
assign n_6407 =  x_1438 & ~n_6334;
assign n_6408 =  i_20 &  n_6334;
assign n_6409 = ~n_6407 & ~n_6408;
assign n_6410 =  x_1438 & ~n_6409;
assign n_6411 = ~x_1438 &  n_6409;
assign n_6412 = ~n_6410 & ~n_6411;
assign n_6413 =  x_1437 & ~n_6334;
assign n_6414 =  i_19 &  n_6334;
assign n_6415 = ~n_6413 & ~n_6414;
assign n_6416 =  x_1437 & ~n_6415;
assign n_6417 = ~x_1437 &  n_6415;
assign n_6418 = ~n_6416 & ~n_6417;
assign n_6419 =  x_1436 & ~n_6334;
assign n_6420 =  i_18 &  n_6334;
assign n_6421 = ~n_6419 & ~n_6420;
assign n_6422 =  x_1436 & ~n_6421;
assign n_6423 = ~x_1436 &  n_6421;
assign n_6424 = ~n_6422 & ~n_6423;
assign n_6425 =  x_1435 & ~n_6334;
assign n_6426 =  i_17 &  n_6334;
assign n_6427 = ~n_6425 & ~n_6426;
assign n_6428 =  x_1435 & ~n_6427;
assign n_6429 = ~x_1435 &  n_6427;
assign n_6430 = ~n_6428 & ~n_6429;
assign n_6431 =  x_1434 & ~n_6334;
assign n_6432 =  i_16 &  n_6334;
assign n_6433 = ~n_6431 & ~n_6432;
assign n_6434 =  x_1434 & ~n_6433;
assign n_6435 = ~x_1434 &  n_6433;
assign n_6436 = ~n_6434 & ~n_6435;
assign n_6437 =  x_1433 & ~n_6334;
assign n_6438 =  i_15 &  n_6334;
assign n_6439 = ~n_6437 & ~n_6438;
assign n_6440 =  x_1433 & ~n_6439;
assign n_6441 = ~x_1433 &  n_6439;
assign n_6442 = ~n_6440 & ~n_6441;
assign n_6443 =  x_1432 & ~n_6334;
assign n_6444 =  i_14 &  n_6334;
assign n_6445 = ~n_6443 & ~n_6444;
assign n_6446 =  x_1432 & ~n_6445;
assign n_6447 = ~x_1432 &  n_6445;
assign n_6448 = ~n_6446 & ~n_6447;
assign n_6449 =  x_1431 & ~n_6334;
assign n_6450 =  i_13 &  n_6334;
assign n_6451 = ~n_6449 & ~n_6450;
assign n_6452 =  x_1431 & ~n_6451;
assign n_6453 = ~x_1431 &  n_6451;
assign n_6454 = ~n_6452 & ~n_6453;
assign n_6455 =  x_1430 & ~n_6334;
assign n_6456 =  i_12 &  n_6334;
assign n_6457 = ~n_6455 & ~n_6456;
assign n_6458 =  x_1430 & ~n_6457;
assign n_6459 = ~x_1430 &  n_6457;
assign n_6460 = ~n_6458 & ~n_6459;
assign n_6461 =  x_1429 & ~n_6334;
assign n_6462 =  i_11 &  n_6334;
assign n_6463 = ~n_6461 & ~n_6462;
assign n_6464 =  x_1429 & ~n_6463;
assign n_6465 = ~x_1429 &  n_6463;
assign n_6466 = ~n_6464 & ~n_6465;
assign n_6467 =  x_1428 & ~n_6334;
assign n_6468 =  i_10 &  n_6334;
assign n_6469 = ~n_6467 & ~n_6468;
assign n_6470 =  x_1428 & ~n_6469;
assign n_6471 = ~x_1428 &  n_6469;
assign n_6472 = ~n_6470 & ~n_6471;
assign n_6473 =  x_1427 & ~n_6334;
assign n_6474 =  i_9 &  n_6334;
assign n_6475 = ~n_6473 & ~n_6474;
assign n_6476 =  x_1427 & ~n_6475;
assign n_6477 = ~x_1427 &  n_6475;
assign n_6478 = ~n_6476 & ~n_6477;
assign n_6479 =  x_1426 & ~n_6334;
assign n_6480 =  i_8 &  n_6334;
assign n_6481 = ~n_6479 & ~n_6480;
assign n_6482 =  x_1426 & ~n_6481;
assign n_6483 = ~x_1426 &  n_6481;
assign n_6484 = ~n_6482 & ~n_6483;
assign n_6485 =  x_1425 & ~n_6334;
assign n_6486 =  i_7 &  n_6334;
assign n_6487 = ~n_6485 & ~n_6486;
assign n_6488 =  x_1425 & ~n_6487;
assign n_6489 = ~x_1425 &  n_6487;
assign n_6490 = ~n_6488 & ~n_6489;
assign n_6491 =  x_1424 & ~n_6334;
assign n_6492 =  i_6 &  n_6334;
assign n_6493 = ~n_6491 & ~n_6492;
assign n_6494 =  x_1424 & ~n_6493;
assign n_6495 = ~x_1424 &  n_6493;
assign n_6496 = ~n_6494 & ~n_6495;
assign n_6497 =  x_1423 & ~n_6334;
assign n_6498 =  i_5 &  n_6334;
assign n_6499 = ~n_6497 & ~n_6498;
assign n_6500 =  x_1423 & ~n_6499;
assign n_6501 = ~x_1423 &  n_6499;
assign n_6502 = ~n_6500 & ~n_6501;
assign n_6503 =  x_1422 & ~n_6334;
assign n_6504 =  i_4 &  n_6334;
assign n_6505 = ~n_6503 & ~n_6504;
assign n_6506 =  x_1422 & ~n_6505;
assign n_6507 = ~x_1422 &  n_6505;
assign n_6508 = ~n_6506 & ~n_6507;
assign n_6509 =  x_1421 & ~n_6334;
assign n_6510 =  i_3 &  n_6334;
assign n_6511 = ~n_6509 & ~n_6510;
assign n_6512 =  x_1421 & ~n_6511;
assign n_6513 = ~x_1421 &  n_6511;
assign n_6514 = ~n_6512 & ~n_6513;
assign n_6515 =  x_1420 & ~n_6334;
assign n_6516 =  i_2 &  n_6334;
assign n_6517 = ~n_6515 & ~n_6516;
assign n_6518 =  x_1420 & ~n_6517;
assign n_6519 = ~x_1420 &  n_6517;
assign n_6520 = ~n_6518 & ~n_6519;
assign n_6521 =  x_1419 & ~n_6334;
assign n_6522 =  i_1 &  n_6334;
assign n_6523 = ~n_6521 & ~n_6522;
assign n_6524 =  x_1419 & ~n_6523;
assign n_6525 = ~x_1419 &  n_6523;
assign n_6526 = ~n_6524 & ~n_6525;
assign n_6527 =  n_389 &  n_1708;
assign n_6528 =  n_386 &  n_6527;
assign n_6529 =  x_41 &  n_6528;
assign n_6530 =  n_2 &  n_3861;
assign n_6531 =  n_6530 &  n_785;
assign n_6532 =  n_388 &  n_2100;
assign n_6533 = ~x_42 &  n_3663;
assign n_6534 =  n_6532 &  n_6533;
assign n_6535 = ~n_6531 & ~n_6534;
assign n_6536 = ~n_6529 &  n_6535;
assign n_6537 =  x_1418 &  n_6536;
assign n_6538 =  x_586 &  x_2154;
assign n_6539 = ~x_586 & ~x_2154;
assign n_6540 = ~n_6538 & ~n_6539;
assign n_6541 =  n_6531 &  n_6540;
assign n_6542 =  x_2250 &  x_2762;
assign n_6543 = ~x_2250 & ~x_2762;
assign n_6544 = ~n_6542 & ~n_6543;
assign n_6545 =  n_6534 &  n_6544;
assign n_6546 = ~n_6541 & ~n_6545;
assign n_6547 = ~n_6537 &  n_6546;
assign n_6548 =  x_1418 & ~n_6547;
assign n_6549 = ~x_1418 &  n_6547;
assign n_6550 = ~n_6548 & ~n_6549;
assign n_6551 =  x_1417 &  n_6536;
assign n_6552 = ~x_2761 & ~x_2762;
assign n_6553 =  x_2761 &  x_2762;
assign n_6554 = ~n_6552 & ~n_6553;
assign n_6555 =  x_2249 &  n_6554;
assign n_6556 = ~x_2249 & ~n_6554;
assign n_6557 = ~n_6555 & ~n_6556;
assign n_6558 =  n_6542 &  n_6557;
assign n_6559 = ~n_6542 & ~n_6557;
assign n_6560 =  n_6534 & ~n_6559;
assign n_6561 = ~n_6558 &  n_6560;
assign n_6562 = ~x_2153 & ~x_2154;
assign n_6563 =  x_2153 &  x_2154;
assign n_6564 = ~n_6562 & ~n_6563;
assign n_6565 =  x_585 &  n_6564;
assign n_6566 = ~x_585 & ~n_6564;
assign n_6567 = ~n_6565 & ~n_6566;
assign n_6568 = ~n_6538 & ~n_6567;
assign n_6569 =  n_6538 &  n_6567;
assign n_6570 =  n_6531 & ~n_6569;
assign n_6571 = ~n_6568 &  n_6570;
assign n_6572 = ~n_6561 & ~n_6571;
assign n_6573 = ~n_6551 &  n_6572;
assign n_6574 =  x_1417 & ~n_6573;
assign n_6575 = ~x_1417 &  n_6573;
assign n_6576 = ~n_6574 & ~n_6575;
assign n_6577 = ~x_2152 &  n_6562;
assign n_6578 =  x_2152 & ~n_6562;
assign n_6579 = ~n_6577 & ~n_6578;
assign n_6580 = ~x_585 &  x_2153;
assign n_6581 =  n_6538 & ~n_6580;
assign n_6582 = ~n_6581 & ~n_6565;
assign n_6583 =  n_6579 & ~n_6582;
assign n_6584 = ~n_6579 &  n_6582;
assign n_6585 = ~n_6583 & ~n_6584;
assign n_6586 = ~x_584 & ~n_6585;
assign n_6587 =  x_584 & ~n_6584;
assign n_6588 = ~n_6583 &  n_6587;
assign n_6589 =  n_6531 & ~n_6588;
assign n_6590 = ~n_6586 &  n_6589;
assign n_6591 =  x_1416 &  n_6536;
assign n_6592 = ~x_2760 &  n_6552;
assign n_6593 =  x_2760 & ~n_6552;
assign n_6594 = ~n_6592 & ~n_6593;
assign n_6595 = ~x_2249 &  x_2761;
assign n_6596 =  n_6542 & ~n_6595;
assign n_6597 = ~n_6596 & ~n_6555;
assign n_6598 =  n_6594 & ~n_6597;
assign n_6599 = ~n_6594 &  n_6597;
assign n_6600 = ~n_6598 & ~n_6599;
assign n_6601 = ~x_2248 & ~n_6600;
assign n_6602 =  x_2248 & ~n_6599;
assign n_6603 = ~n_6598 &  n_6602;
assign n_6604 =  n_6534 & ~n_6603;
assign n_6605 = ~n_6601 &  n_6604;
assign n_6606 = ~n_6591 & ~n_6605;
assign n_6607 = ~n_6590 &  n_6606;
assign n_6608 =  x_1416 & ~n_6607;
assign n_6609 = ~x_1416 &  n_6607;
assign n_6610 = ~n_6608 & ~n_6609;
assign n_6611 = ~x_2151 &  n_6577;
assign n_6612 =  x_2151 & ~n_6577;
assign n_6613 = ~n_6611 & ~n_6612;
assign n_6614 = ~n_6583 & ~n_6587;
assign n_6615 =  n_6613 & ~n_6614;
assign n_6616 = ~n_6613 &  n_6614;
assign n_6617 = ~n_6615 & ~n_6616;
assign n_6618 = ~x_583 & ~n_6617;
assign n_6619 =  x_583 & ~n_6616;
assign n_6620 = ~n_6615 &  n_6619;
assign n_6621 =  n_6531 & ~n_6620;
assign n_6622 = ~n_6618 &  n_6621;
assign n_6623 =  x_1415 &  n_6536;
assign n_6624 = ~x_2759 &  n_6592;
assign n_6625 =  x_2759 & ~n_6592;
assign n_6626 = ~n_6624 & ~n_6625;
assign n_6627 = ~n_6598 & ~n_6602;
assign n_6628 =  n_6626 & ~n_6627;
assign n_6629 = ~n_6626 &  n_6627;
assign n_6630 = ~n_6628 & ~n_6629;
assign n_6631 = ~x_2247 & ~n_6630;
assign n_6632 =  x_2247 & ~n_6629;
assign n_6633 = ~n_6628 &  n_6632;
assign n_6634 =  n_6534 & ~n_6633;
assign n_6635 = ~n_6631 &  n_6634;
assign n_6636 = ~n_6623 & ~n_6635;
assign n_6637 = ~n_6622 &  n_6636;
assign n_6638 =  x_1415 & ~n_6637;
assign n_6639 = ~x_1415 &  n_6637;
assign n_6640 = ~n_6638 & ~n_6639;
assign n_6641 = ~x_2758 &  n_6624;
assign n_6642 =  x_2758 & ~n_6624;
assign n_6643 = ~n_6641 & ~n_6642;
assign n_6644 = ~n_6628 & ~n_6632;
assign n_6645 =  n_6643 & ~n_6644;
assign n_6646 = ~n_6643 &  n_6644;
assign n_6647 = ~n_6645 & ~n_6646;
assign n_6648 = ~x_2246 & ~n_6647;
assign n_6649 =  x_2246 & ~n_6646;
assign n_6650 = ~n_6645 &  n_6649;
assign n_6651 =  n_6534 & ~n_6650;
assign n_6652 = ~n_6648 &  n_6651;
assign n_6653 =  x_1414 &  n_6536;
assign n_6654 = ~x_2150 &  n_6611;
assign n_6655 =  x_2150 & ~n_6611;
assign n_6656 = ~n_6654 & ~n_6655;
assign n_6657 = ~n_6615 & ~n_6619;
assign n_6658 =  n_6656 & ~n_6657;
assign n_6659 = ~n_6656 &  n_6657;
assign n_6660 = ~n_6658 & ~n_6659;
assign n_6661 = ~x_582 & ~n_6660;
assign n_6662 =  x_582 & ~n_6659;
assign n_6663 = ~n_6658 &  n_6662;
assign n_6664 =  n_6531 & ~n_6663;
assign n_6665 = ~n_6661 &  n_6664;
assign n_6666 = ~n_6653 & ~n_6665;
assign n_6667 = ~n_6652 &  n_6666;
assign n_6668 =  x_1414 & ~n_6667;
assign n_6669 = ~x_1414 &  n_6667;
assign n_6670 = ~n_6668 & ~n_6669;
assign n_6671 = ~x_2757 &  n_6641;
assign n_6672 =  x_2757 & ~n_6641;
assign n_6673 = ~n_6671 & ~n_6672;
assign n_6674 = ~n_6645 & ~n_6649;
assign n_6675 =  n_6673 & ~n_6674;
assign n_6676 = ~n_6673 &  n_6674;
assign n_6677 = ~n_6675 & ~n_6676;
assign n_6678 = ~x_2245 & ~n_6677;
assign n_6679 =  x_2245 & ~n_6676;
assign n_6680 = ~n_6675 &  n_6679;
assign n_6681 =  n_6534 & ~n_6680;
assign n_6682 = ~n_6678 &  n_6681;
assign n_6683 =  x_1413 &  n_6536;
assign n_6684 = ~x_2149 &  n_6654;
assign n_6685 =  x_2149 & ~n_6654;
assign n_6686 = ~n_6684 & ~n_6685;
assign n_6687 = ~n_6658 & ~n_6662;
assign n_6688 =  n_6686 & ~n_6687;
assign n_6689 = ~n_6686 &  n_6687;
assign n_6690 = ~n_6688 & ~n_6689;
assign n_6691 = ~x_581 & ~n_6690;
assign n_6692 =  x_581 & ~n_6689;
assign n_6693 = ~n_6688 &  n_6692;
assign n_6694 =  n_6531 & ~n_6693;
assign n_6695 = ~n_6691 &  n_6694;
assign n_6696 = ~n_6683 & ~n_6695;
assign n_6697 = ~n_6682 &  n_6696;
assign n_6698 =  x_1413 & ~n_6697;
assign n_6699 = ~x_1413 &  n_6697;
assign n_6700 = ~n_6698 & ~n_6699;
assign n_6701 = ~x_2756 &  n_6671;
assign n_6702 =  x_2756 & ~n_6671;
assign n_6703 = ~n_6701 & ~n_6702;
assign n_6704 = ~n_6675 & ~n_6679;
assign n_6705 =  n_6703 & ~n_6704;
assign n_6706 = ~n_6703 &  n_6704;
assign n_6707 = ~n_6705 & ~n_6706;
assign n_6708 = ~x_2244 & ~n_6707;
assign n_6709 =  x_2244 & ~n_6706;
assign n_6710 = ~n_6705 &  n_6709;
assign n_6711 =  n_6534 & ~n_6710;
assign n_6712 = ~n_6708 &  n_6711;
assign n_6713 =  x_1412 &  n_6536;
assign n_6714 = ~x_2148 &  n_6684;
assign n_6715 =  x_2148 & ~n_6684;
assign n_6716 = ~n_6714 & ~n_6715;
assign n_6717 = ~n_6688 & ~n_6692;
assign n_6718 =  n_6716 & ~n_6717;
assign n_6719 = ~n_6716 &  n_6717;
assign n_6720 = ~n_6718 & ~n_6719;
assign n_6721 = ~x_580 & ~n_6720;
assign n_6722 =  x_580 & ~n_6719;
assign n_6723 = ~n_6718 &  n_6722;
assign n_6724 =  n_6531 & ~n_6723;
assign n_6725 = ~n_6721 &  n_6724;
assign n_6726 = ~n_6713 & ~n_6725;
assign n_6727 = ~n_6712 &  n_6726;
assign n_6728 =  x_1412 & ~n_6727;
assign n_6729 = ~x_1412 &  n_6727;
assign n_6730 = ~n_6728 & ~n_6729;
assign n_6731 = ~x_2755 &  n_6701;
assign n_6732 =  x_2755 & ~n_6701;
assign n_6733 = ~n_6731 & ~n_6732;
assign n_6734 = ~n_6705 & ~n_6709;
assign n_6735 =  n_6733 & ~n_6734;
assign n_6736 = ~n_6733 &  n_6734;
assign n_6737 = ~n_6735 & ~n_6736;
assign n_6738 = ~x_2243 & ~n_6737;
assign n_6739 =  x_2243 & ~n_6736;
assign n_6740 = ~n_6735 &  n_6739;
assign n_6741 =  n_6534 & ~n_6740;
assign n_6742 = ~n_6738 &  n_6741;
assign n_6743 =  x_1411 &  n_6536;
assign n_6744 = ~x_2147 &  n_6714;
assign n_6745 =  x_2147 & ~n_6714;
assign n_6746 = ~n_6744 & ~n_6745;
assign n_6747 = ~n_6718 & ~n_6722;
assign n_6748 =  n_6746 & ~n_6747;
assign n_6749 = ~n_6746 &  n_6747;
assign n_6750 = ~n_6748 & ~n_6749;
assign n_6751 = ~x_579 & ~n_6750;
assign n_6752 =  x_579 & ~n_6749;
assign n_6753 = ~n_6748 &  n_6752;
assign n_6754 =  n_6531 & ~n_6753;
assign n_6755 = ~n_6751 &  n_6754;
assign n_6756 = ~n_6743 & ~n_6755;
assign n_6757 = ~n_6742 &  n_6756;
assign n_6758 =  x_1411 & ~n_6757;
assign n_6759 = ~x_1411 &  n_6757;
assign n_6760 = ~n_6758 & ~n_6759;
assign n_6761 = ~x_2754 &  n_6731;
assign n_6762 =  x_2754 & ~n_6731;
assign n_6763 = ~n_6761 & ~n_6762;
assign n_6764 = ~n_6735 & ~n_6739;
assign n_6765 =  n_6763 & ~n_6764;
assign n_6766 = ~n_6763 &  n_6764;
assign n_6767 = ~n_6765 & ~n_6766;
assign n_6768 = ~x_2242 & ~n_6767;
assign n_6769 =  x_2242 & ~n_6766;
assign n_6770 = ~n_6765 &  n_6769;
assign n_6771 =  n_6534 & ~n_6770;
assign n_6772 = ~n_6768 &  n_6771;
assign n_6773 =  x_1410 &  n_6536;
assign n_6774 = ~x_2146 &  n_6744;
assign n_6775 =  x_2146 & ~n_6744;
assign n_6776 = ~n_6774 & ~n_6775;
assign n_6777 = ~n_6748 & ~n_6752;
assign n_6778 =  n_6776 & ~n_6777;
assign n_6779 = ~n_6776 &  n_6777;
assign n_6780 = ~n_6778 & ~n_6779;
assign n_6781 = ~x_578 & ~n_6780;
assign n_6782 =  x_578 & ~n_6779;
assign n_6783 = ~n_6778 &  n_6782;
assign n_6784 =  n_6531 & ~n_6783;
assign n_6785 = ~n_6781 &  n_6784;
assign n_6786 = ~n_6773 & ~n_6785;
assign n_6787 = ~n_6772 &  n_6786;
assign n_6788 =  x_1410 & ~n_6787;
assign n_6789 = ~x_1410 &  n_6787;
assign n_6790 = ~n_6788 & ~n_6789;
assign n_6791 = ~x_2753 &  n_6761;
assign n_6792 =  x_2753 & ~n_6761;
assign n_6793 = ~n_6791 & ~n_6792;
assign n_6794 = ~n_6765 & ~n_6769;
assign n_6795 =  n_6793 & ~n_6794;
assign n_6796 = ~n_6793 &  n_6794;
assign n_6797 = ~n_6795 & ~n_6796;
assign n_6798 = ~x_2241 & ~n_6797;
assign n_6799 =  x_2241 & ~n_6796;
assign n_6800 = ~n_6795 &  n_6799;
assign n_6801 =  n_6534 & ~n_6800;
assign n_6802 = ~n_6798 &  n_6801;
assign n_6803 =  x_1409 &  n_6536;
assign n_6804 = ~x_2145 &  n_6774;
assign n_6805 =  x_2145 & ~n_6774;
assign n_6806 = ~n_6804 & ~n_6805;
assign n_6807 = ~n_6778 & ~n_6782;
assign n_6808 =  n_6806 & ~n_6807;
assign n_6809 = ~n_6806 &  n_6807;
assign n_6810 = ~n_6808 & ~n_6809;
assign n_6811 = ~x_577 & ~n_6810;
assign n_6812 =  x_577 & ~n_6809;
assign n_6813 = ~n_6808 &  n_6812;
assign n_6814 =  n_6531 & ~n_6813;
assign n_6815 = ~n_6811 &  n_6814;
assign n_6816 = ~n_6803 & ~n_6815;
assign n_6817 = ~n_6802 &  n_6816;
assign n_6818 =  x_1409 & ~n_6817;
assign n_6819 = ~x_1409 &  n_6817;
assign n_6820 = ~n_6818 & ~n_6819;
assign n_6821 = ~x_2752 &  n_6791;
assign n_6822 =  x_2752 & ~n_6791;
assign n_6823 = ~n_6821 & ~n_6822;
assign n_6824 = ~n_6795 & ~n_6799;
assign n_6825 =  n_6823 & ~n_6824;
assign n_6826 = ~n_6823 &  n_6824;
assign n_6827 = ~n_6825 & ~n_6826;
assign n_6828 = ~x_2240 & ~n_6827;
assign n_6829 =  x_2240 & ~n_6826;
assign n_6830 = ~n_6825 &  n_6829;
assign n_6831 =  n_6534 & ~n_6830;
assign n_6832 = ~n_6828 &  n_6831;
assign n_6833 =  x_1408 &  n_6536;
assign n_6834 = ~x_2144 &  n_6804;
assign n_6835 =  x_2144 & ~n_6804;
assign n_6836 = ~n_6834 & ~n_6835;
assign n_6837 = ~n_6808 & ~n_6812;
assign n_6838 =  n_6836 & ~n_6837;
assign n_6839 = ~n_6836 &  n_6837;
assign n_6840 = ~n_6838 & ~n_6839;
assign n_6841 = ~x_576 & ~n_6840;
assign n_6842 =  x_576 & ~n_6839;
assign n_6843 = ~n_6838 &  n_6842;
assign n_6844 =  n_6531 & ~n_6843;
assign n_6845 = ~n_6841 &  n_6844;
assign n_6846 = ~n_6833 & ~n_6845;
assign n_6847 = ~n_6832 &  n_6846;
assign n_6848 =  x_1408 & ~n_6847;
assign n_6849 = ~x_1408 &  n_6847;
assign n_6850 = ~n_6848 & ~n_6849;
assign n_6851 = ~x_2751 &  n_6821;
assign n_6852 =  x_2751 & ~n_6821;
assign n_6853 = ~n_6851 & ~n_6852;
assign n_6854 = ~n_6825 & ~n_6829;
assign n_6855 =  n_6853 & ~n_6854;
assign n_6856 = ~n_6853 &  n_6854;
assign n_6857 = ~n_6855 & ~n_6856;
assign n_6858 = ~x_2239 & ~n_6857;
assign n_6859 =  x_2239 & ~n_6856;
assign n_6860 = ~n_6855 &  n_6859;
assign n_6861 =  n_6534 & ~n_6860;
assign n_6862 = ~n_6858 &  n_6861;
assign n_6863 =  x_1407 &  n_6536;
assign n_6864 = ~x_2143 &  n_6834;
assign n_6865 =  x_2143 & ~n_6834;
assign n_6866 = ~n_6864 & ~n_6865;
assign n_6867 = ~n_6838 & ~n_6842;
assign n_6868 =  n_6866 & ~n_6867;
assign n_6869 = ~n_6866 &  n_6867;
assign n_6870 = ~n_6868 & ~n_6869;
assign n_6871 = ~x_575 & ~n_6870;
assign n_6872 =  x_575 & ~n_6869;
assign n_6873 = ~n_6868 &  n_6872;
assign n_6874 =  n_6531 & ~n_6873;
assign n_6875 = ~n_6871 &  n_6874;
assign n_6876 = ~n_6863 & ~n_6875;
assign n_6877 = ~n_6862 &  n_6876;
assign n_6878 =  x_1407 & ~n_6877;
assign n_6879 = ~x_1407 &  n_6877;
assign n_6880 = ~n_6878 & ~n_6879;
assign n_6881 = ~x_2750 &  n_6851;
assign n_6882 =  x_2750 & ~n_6851;
assign n_6883 = ~n_6881 & ~n_6882;
assign n_6884 = ~n_6855 & ~n_6859;
assign n_6885 =  n_6883 & ~n_6884;
assign n_6886 = ~n_6883 &  n_6884;
assign n_6887 = ~n_6885 & ~n_6886;
assign n_6888 = ~x_2238 & ~n_6887;
assign n_6889 =  x_2238 & ~n_6886;
assign n_6890 = ~n_6885 &  n_6889;
assign n_6891 =  n_6534 & ~n_6890;
assign n_6892 = ~n_6888 &  n_6891;
assign n_6893 =  x_1406 &  n_6536;
assign n_6894 = ~x_2142 &  n_6864;
assign n_6895 =  x_2142 & ~n_6864;
assign n_6896 = ~n_6894 & ~n_6895;
assign n_6897 = ~n_6868 & ~n_6872;
assign n_6898 =  n_6896 & ~n_6897;
assign n_6899 = ~n_6896 &  n_6897;
assign n_6900 = ~n_6898 & ~n_6899;
assign n_6901 = ~x_574 & ~n_6900;
assign n_6902 =  x_574 & ~n_6899;
assign n_6903 = ~n_6898 &  n_6902;
assign n_6904 =  n_6531 & ~n_6903;
assign n_6905 = ~n_6901 &  n_6904;
assign n_6906 = ~n_6893 & ~n_6905;
assign n_6907 = ~n_6892 &  n_6906;
assign n_6908 =  x_1406 & ~n_6907;
assign n_6909 = ~x_1406 &  n_6907;
assign n_6910 = ~n_6908 & ~n_6909;
assign n_6911 = ~x_2749 &  n_6881;
assign n_6912 =  x_2749 & ~n_6881;
assign n_6913 = ~n_6911 & ~n_6912;
assign n_6914 = ~n_6885 & ~n_6889;
assign n_6915 =  n_6913 & ~n_6914;
assign n_6916 = ~n_6913 &  n_6914;
assign n_6917 = ~n_6915 & ~n_6916;
assign n_6918 = ~x_2237 & ~n_6917;
assign n_6919 =  x_2237 & ~n_6916;
assign n_6920 = ~n_6915 &  n_6919;
assign n_6921 =  n_6534 & ~n_6920;
assign n_6922 = ~n_6918 &  n_6921;
assign n_6923 =  x_1405 &  n_6536;
assign n_6924 = ~x_2141 &  n_6894;
assign n_6925 =  x_2141 & ~n_6894;
assign n_6926 = ~n_6924 & ~n_6925;
assign n_6927 = ~n_6898 & ~n_6902;
assign n_6928 =  n_6926 & ~n_6927;
assign n_6929 = ~n_6926 &  n_6927;
assign n_6930 = ~n_6928 & ~n_6929;
assign n_6931 = ~x_573 & ~n_6930;
assign n_6932 =  x_573 & ~n_6929;
assign n_6933 = ~n_6928 &  n_6932;
assign n_6934 =  n_6531 & ~n_6933;
assign n_6935 = ~n_6931 &  n_6934;
assign n_6936 = ~n_6923 & ~n_6935;
assign n_6937 = ~n_6922 &  n_6936;
assign n_6938 =  x_1405 & ~n_6937;
assign n_6939 = ~x_1405 &  n_6937;
assign n_6940 = ~n_6938 & ~n_6939;
assign n_6941 = ~x_2748 &  n_6911;
assign n_6942 =  x_2748 & ~n_6911;
assign n_6943 = ~n_6941 & ~n_6942;
assign n_6944 = ~n_6915 & ~n_6919;
assign n_6945 =  n_6943 & ~n_6944;
assign n_6946 = ~n_6943 &  n_6944;
assign n_6947 = ~n_6945 & ~n_6946;
assign n_6948 = ~x_2236 & ~n_6947;
assign n_6949 =  x_2236 & ~n_6946;
assign n_6950 = ~n_6945 &  n_6949;
assign n_6951 =  n_6534 & ~n_6950;
assign n_6952 = ~n_6948 &  n_6951;
assign n_6953 =  x_1404 &  n_6536;
assign n_6954 = ~x_2140 &  n_6924;
assign n_6955 =  x_2140 & ~n_6924;
assign n_6956 = ~n_6954 & ~n_6955;
assign n_6957 = ~n_6928 & ~n_6932;
assign n_6958 =  n_6956 & ~n_6957;
assign n_6959 = ~n_6956 &  n_6957;
assign n_6960 = ~n_6958 & ~n_6959;
assign n_6961 = ~x_572 & ~n_6960;
assign n_6962 =  x_572 & ~n_6959;
assign n_6963 = ~n_6958 &  n_6962;
assign n_6964 =  n_6531 & ~n_6963;
assign n_6965 = ~n_6961 &  n_6964;
assign n_6966 = ~n_6953 & ~n_6965;
assign n_6967 = ~n_6952 &  n_6966;
assign n_6968 =  x_1404 & ~n_6967;
assign n_6969 = ~x_1404 &  n_6967;
assign n_6970 = ~n_6968 & ~n_6969;
assign n_6971 = ~x_2747 &  n_6941;
assign n_6972 =  x_2747 & ~n_6941;
assign n_6973 = ~n_6971 & ~n_6972;
assign n_6974 = ~n_6945 & ~n_6949;
assign n_6975 =  n_6973 & ~n_6974;
assign n_6976 = ~n_6973 &  n_6974;
assign n_6977 = ~n_6975 & ~n_6976;
assign n_6978 = ~x_2235 & ~n_6977;
assign n_6979 =  x_2235 & ~n_6976;
assign n_6980 = ~n_6975 &  n_6979;
assign n_6981 =  n_6534 & ~n_6980;
assign n_6982 = ~n_6978 &  n_6981;
assign n_6983 =  x_1403 &  n_6536;
assign n_6984 = ~x_2139 &  n_6954;
assign n_6985 =  x_2139 & ~n_6954;
assign n_6986 = ~n_6984 & ~n_6985;
assign n_6987 = ~n_6958 & ~n_6962;
assign n_6988 =  n_6986 & ~n_6987;
assign n_6989 = ~n_6986 &  n_6987;
assign n_6990 = ~n_6988 & ~n_6989;
assign n_6991 = ~x_571 & ~n_6990;
assign n_6992 =  x_571 & ~n_6989;
assign n_6993 = ~n_6988 &  n_6992;
assign n_6994 =  n_6531 & ~n_6993;
assign n_6995 = ~n_6991 &  n_6994;
assign n_6996 = ~n_6983 & ~n_6995;
assign n_6997 = ~n_6982 &  n_6996;
assign n_6998 =  x_1403 & ~n_6997;
assign n_6999 = ~x_1403 &  n_6997;
assign n_7000 = ~n_6998 & ~n_6999;
assign n_7001 = ~x_2746 &  n_6971;
assign n_7002 =  x_2746 & ~n_6971;
assign n_7003 = ~n_7001 & ~n_7002;
assign n_7004 = ~n_6975 & ~n_6979;
assign n_7005 =  n_7003 & ~n_7004;
assign n_7006 = ~n_7003 &  n_7004;
assign n_7007 = ~n_7005 & ~n_7006;
assign n_7008 = ~x_2234 & ~n_7007;
assign n_7009 =  x_2234 & ~n_7006;
assign n_7010 = ~n_7005 &  n_7009;
assign n_7011 =  n_6534 & ~n_7010;
assign n_7012 = ~n_7008 &  n_7011;
assign n_7013 =  x_1402 &  n_6536;
assign n_7014 = ~x_2138 &  n_6984;
assign n_7015 =  x_2138 & ~n_6984;
assign n_7016 = ~n_7014 & ~n_7015;
assign n_7017 = ~n_6988 & ~n_6992;
assign n_7018 =  n_7016 & ~n_7017;
assign n_7019 = ~n_7016 &  n_7017;
assign n_7020 = ~n_7018 & ~n_7019;
assign n_7021 = ~x_570 & ~n_7020;
assign n_7022 =  x_570 & ~n_7019;
assign n_7023 = ~n_7018 &  n_7022;
assign n_7024 =  n_6531 & ~n_7023;
assign n_7025 = ~n_7021 &  n_7024;
assign n_7026 = ~n_7013 & ~n_7025;
assign n_7027 = ~n_7012 &  n_7026;
assign n_7028 =  x_1402 & ~n_7027;
assign n_7029 = ~x_1402 &  n_7027;
assign n_7030 = ~n_7028 & ~n_7029;
assign n_7031 = ~x_2745 &  n_7001;
assign n_7032 =  x_2745 & ~n_7001;
assign n_7033 = ~n_7031 & ~n_7032;
assign n_7034 = ~n_7005 & ~n_7009;
assign n_7035 =  n_7033 & ~n_7034;
assign n_7036 = ~n_7033 &  n_7034;
assign n_7037 = ~n_7035 & ~n_7036;
assign n_7038 = ~x_2233 & ~n_7037;
assign n_7039 =  x_2233 & ~n_7036;
assign n_7040 = ~n_7035 &  n_7039;
assign n_7041 =  n_6534 & ~n_7040;
assign n_7042 = ~n_7038 &  n_7041;
assign n_7043 =  x_1401 &  n_6536;
assign n_7044 = ~x_2137 &  n_7014;
assign n_7045 =  x_2137 & ~n_7014;
assign n_7046 = ~n_7044 & ~n_7045;
assign n_7047 = ~n_7018 & ~n_7022;
assign n_7048 =  n_7046 & ~n_7047;
assign n_7049 = ~n_7046 &  n_7047;
assign n_7050 = ~n_7048 & ~n_7049;
assign n_7051 = ~x_569 & ~n_7050;
assign n_7052 =  x_569 & ~n_7049;
assign n_7053 = ~n_7048 &  n_7052;
assign n_7054 =  n_6531 & ~n_7053;
assign n_7055 = ~n_7051 &  n_7054;
assign n_7056 = ~n_7043 & ~n_7055;
assign n_7057 = ~n_7042 &  n_7056;
assign n_7058 =  x_1401 & ~n_7057;
assign n_7059 = ~x_1401 &  n_7057;
assign n_7060 = ~n_7058 & ~n_7059;
assign n_7061 = ~x_2744 &  n_7031;
assign n_7062 =  x_2744 & ~n_7031;
assign n_7063 = ~n_7061 & ~n_7062;
assign n_7064 = ~n_7035 & ~n_7039;
assign n_7065 =  n_7063 & ~n_7064;
assign n_7066 = ~n_7063 &  n_7064;
assign n_7067 = ~n_7065 & ~n_7066;
assign n_7068 = ~x_2232 & ~n_7067;
assign n_7069 =  x_2232 & ~n_7066;
assign n_7070 = ~n_7065 &  n_7069;
assign n_7071 =  n_6534 & ~n_7070;
assign n_7072 = ~n_7068 &  n_7071;
assign n_7073 =  x_1400 &  n_6536;
assign n_7074 = ~x_2136 &  n_7044;
assign n_7075 =  x_2136 & ~n_7044;
assign n_7076 = ~n_7074 & ~n_7075;
assign n_7077 = ~n_7048 & ~n_7052;
assign n_7078 =  n_7076 & ~n_7077;
assign n_7079 = ~n_7076 &  n_7077;
assign n_7080 = ~n_7078 & ~n_7079;
assign n_7081 = ~x_568 & ~n_7080;
assign n_7082 =  x_568 & ~n_7079;
assign n_7083 = ~n_7078 &  n_7082;
assign n_7084 =  n_6531 & ~n_7083;
assign n_7085 = ~n_7081 &  n_7084;
assign n_7086 = ~n_7073 & ~n_7085;
assign n_7087 = ~n_7072 &  n_7086;
assign n_7088 =  x_1400 & ~n_7087;
assign n_7089 = ~x_1400 &  n_7087;
assign n_7090 = ~n_7088 & ~n_7089;
assign n_7091 = ~x_2743 &  n_7061;
assign n_7092 =  x_2743 & ~n_7061;
assign n_7093 = ~n_7091 & ~n_7092;
assign n_7094 = ~n_7065 & ~n_7069;
assign n_7095 =  n_7093 & ~n_7094;
assign n_7096 = ~n_7093 &  n_7094;
assign n_7097 = ~n_7095 & ~n_7096;
assign n_7098 = ~x_2231 & ~n_7097;
assign n_7099 =  x_2231 & ~n_7096;
assign n_7100 = ~n_7095 &  n_7099;
assign n_7101 =  n_6534 & ~n_7100;
assign n_7102 = ~n_7098 &  n_7101;
assign n_7103 =  x_1399 &  n_6536;
assign n_7104 = ~x_2135 &  n_7074;
assign n_7105 =  x_2135 & ~n_7074;
assign n_7106 = ~n_7104 & ~n_7105;
assign n_7107 = ~n_7078 & ~n_7082;
assign n_7108 =  n_7106 & ~n_7107;
assign n_7109 = ~n_7106 &  n_7107;
assign n_7110 = ~n_7108 & ~n_7109;
assign n_7111 = ~x_567 & ~n_7110;
assign n_7112 =  x_567 & ~n_7109;
assign n_7113 = ~n_7108 &  n_7112;
assign n_7114 =  n_6531 & ~n_7113;
assign n_7115 = ~n_7111 &  n_7114;
assign n_7116 = ~n_7103 & ~n_7115;
assign n_7117 = ~n_7102 &  n_7116;
assign n_7118 =  x_1399 & ~n_7117;
assign n_7119 = ~x_1399 &  n_7117;
assign n_7120 = ~n_7118 & ~n_7119;
assign n_7121 = ~x_2742 &  n_7091;
assign n_7122 =  x_2742 & ~n_7091;
assign n_7123 = ~n_7121 & ~n_7122;
assign n_7124 = ~n_7095 & ~n_7099;
assign n_7125 =  n_7123 & ~n_7124;
assign n_7126 = ~n_7123 &  n_7124;
assign n_7127 = ~n_7125 & ~n_7126;
assign n_7128 = ~x_2230 & ~n_7127;
assign n_7129 =  x_2230 & ~n_7126;
assign n_7130 = ~n_7125 &  n_7129;
assign n_7131 =  n_6534 & ~n_7130;
assign n_7132 = ~n_7128 &  n_7131;
assign n_7133 =  x_1398 &  n_6536;
assign n_7134 = ~x_2134 &  n_7104;
assign n_7135 =  x_2134 & ~n_7104;
assign n_7136 = ~n_7134 & ~n_7135;
assign n_7137 = ~n_7108 & ~n_7112;
assign n_7138 =  n_7136 & ~n_7137;
assign n_7139 = ~n_7136 &  n_7137;
assign n_7140 = ~n_7138 & ~n_7139;
assign n_7141 = ~x_566 & ~n_7140;
assign n_7142 =  x_566 & ~n_7139;
assign n_7143 = ~n_7138 &  n_7142;
assign n_7144 =  n_6531 & ~n_7143;
assign n_7145 = ~n_7141 &  n_7144;
assign n_7146 = ~n_7133 & ~n_7145;
assign n_7147 = ~n_7132 &  n_7146;
assign n_7148 =  x_1398 & ~n_7147;
assign n_7149 = ~x_1398 &  n_7147;
assign n_7150 = ~n_7148 & ~n_7149;
assign n_7151 = ~x_2741 &  n_7121;
assign n_7152 =  x_2741 & ~n_7121;
assign n_7153 = ~n_7151 & ~n_7152;
assign n_7154 = ~n_7125 & ~n_7129;
assign n_7155 =  n_7153 & ~n_7154;
assign n_7156 = ~n_7153 &  n_7154;
assign n_7157 = ~n_7155 & ~n_7156;
assign n_7158 = ~x_2229 & ~n_7157;
assign n_7159 =  x_2229 & ~n_7156;
assign n_7160 = ~n_7155 &  n_7159;
assign n_7161 =  n_6534 & ~n_7160;
assign n_7162 = ~n_7158 &  n_7161;
assign n_7163 =  x_1397 &  n_6536;
assign n_7164 = ~x_2133 &  n_7134;
assign n_7165 =  x_2133 & ~n_7134;
assign n_7166 = ~n_7164 & ~n_7165;
assign n_7167 = ~n_7138 & ~n_7142;
assign n_7168 =  n_7166 & ~n_7167;
assign n_7169 = ~n_7166 &  n_7167;
assign n_7170 = ~n_7168 & ~n_7169;
assign n_7171 = ~x_565 & ~n_7170;
assign n_7172 =  x_565 & ~n_7169;
assign n_7173 = ~n_7168 &  n_7172;
assign n_7174 =  n_6531 & ~n_7173;
assign n_7175 = ~n_7171 &  n_7174;
assign n_7176 = ~n_7163 & ~n_7175;
assign n_7177 = ~n_7162 &  n_7176;
assign n_7178 =  x_1397 & ~n_7177;
assign n_7179 = ~x_1397 &  n_7177;
assign n_7180 = ~n_7178 & ~n_7179;
assign n_7181 = ~x_2740 &  n_7151;
assign n_7182 =  x_2740 & ~n_7151;
assign n_7183 = ~n_7181 & ~n_7182;
assign n_7184 = ~n_7155 & ~n_7159;
assign n_7185 =  n_7183 & ~n_7184;
assign n_7186 = ~n_7183 &  n_7184;
assign n_7187 = ~n_7185 & ~n_7186;
assign n_7188 = ~x_2228 & ~n_7187;
assign n_7189 =  x_2228 & ~n_7186;
assign n_7190 = ~n_7185 &  n_7189;
assign n_7191 =  n_6534 & ~n_7190;
assign n_7192 = ~n_7188 &  n_7191;
assign n_7193 =  x_1396 &  n_6536;
assign n_7194 = ~x_2132 &  n_7164;
assign n_7195 =  x_2132 & ~n_7164;
assign n_7196 = ~n_7194 & ~n_7195;
assign n_7197 = ~n_7168 & ~n_7172;
assign n_7198 =  n_7196 & ~n_7197;
assign n_7199 = ~n_7196 &  n_7197;
assign n_7200 = ~n_7198 & ~n_7199;
assign n_7201 = ~x_564 & ~n_7200;
assign n_7202 =  x_564 & ~n_7199;
assign n_7203 = ~n_7198 &  n_7202;
assign n_7204 =  n_6531 & ~n_7203;
assign n_7205 = ~n_7201 &  n_7204;
assign n_7206 = ~n_7193 & ~n_7205;
assign n_7207 = ~n_7192 &  n_7206;
assign n_7208 =  x_1396 & ~n_7207;
assign n_7209 = ~x_1396 &  n_7207;
assign n_7210 = ~n_7208 & ~n_7209;
assign n_7211 = ~x_2739 &  n_7181;
assign n_7212 =  x_2739 & ~n_7181;
assign n_7213 = ~n_7211 & ~n_7212;
assign n_7214 = ~n_7185 & ~n_7189;
assign n_7215 =  n_7213 & ~n_7214;
assign n_7216 = ~n_7213 &  n_7214;
assign n_7217 = ~n_7215 & ~n_7216;
assign n_7218 = ~x_2227 & ~n_7217;
assign n_7219 =  x_2227 & ~n_7216;
assign n_7220 = ~n_7215 &  n_7219;
assign n_7221 =  n_6534 & ~n_7220;
assign n_7222 = ~n_7218 &  n_7221;
assign n_7223 =  x_1395 &  n_6536;
assign n_7224 = ~x_2131 &  n_7194;
assign n_7225 =  x_2131 & ~n_7194;
assign n_7226 = ~n_7224 & ~n_7225;
assign n_7227 = ~n_7198 & ~n_7202;
assign n_7228 =  n_7226 & ~n_7227;
assign n_7229 = ~n_7226 &  n_7227;
assign n_7230 = ~n_7228 & ~n_7229;
assign n_7231 = ~x_563 & ~n_7230;
assign n_7232 =  x_563 & ~n_7229;
assign n_7233 = ~n_7228 &  n_7232;
assign n_7234 =  n_6531 & ~n_7233;
assign n_7235 = ~n_7231 &  n_7234;
assign n_7236 = ~n_7223 & ~n_7235;
assign n_7237 = ~n_7222 &  n_7236;
assign n_7238 =  x_1395 & ~n_7237;
assign n_7239 = ~x_1395 &  n_7237;
assign n_7240 = ~n_7238 & ~n_7239;
assign n_7241 = ~x_2738 &  n_7211;
assign n_7242 =  x_2738 & ~n_7211;
assign n_7243 = ~n_7241 & ~n_7242;
assign n_7244 = ~n_7215 & ~n_7219;
assign n_7245 =  n_7243 & ~n_7244;
assign n_7246 = ~n_7243 &  n_7244;
assign n_7247 = ~n_7245 & ~n_7246;
assign n_7248 = ~x_2226 & ~n_7247;
assign n_7249 =  x_2226 & ~n_7246;
assign n_7250 = ~n_7245 &  n_7249;
assign n_7251 =  n_6534 & ~n_7250;
assign n_7252 = ~n_7248 &  n_7251;
assign n_7253 =  x_1394 &  n_6536;
assign n_7254 = ~x_2130 &  n_7224;
assign n_7255 =  x_2130 & ~n_7224;
assign n_7256 = ~n_7254 & ~n_7255;
assign n_7257 = ~n_7228 & ~n_7232;
assign n_7258 =  n_7256 & ~n_7257;
assign n_7259 = ~n_7256 &  n_7257;
assign n_7260 = ~n_7258 & ~n_7259;
assign n_7261 = ~x_562 & ~n_7260;
assign n_7262 =  x_562 & ~n_7259;
assign n_7263 = ~n_7258 &  n_7262;
assign n_7264 =  n_6531 & ~n_7263;
assign n_7265 = ~n_7261 &  n_7264;
assign n_7266 = ~n_7253 & ~n_7265;
assign n_7267 = ~n_7252 &  n_7266;
assign n_7268 =  x_1394 & ~n_7267;
assign n_7269 = ~x_1394 &  n_7267;
assign n_7270 = ~n_7268 & ~n_7269;
assign n_7271 = ~x_2737 &  n_7241;
assign n_7272 =  x_2737 & ~n_7241;
assign n_7273 = ~n_7271 & ~n_7272;
assign n_7274 = ~n_7245 & ~n_7249;
assign n_7275 =  n_7273 & ~n_7274;
assign n_7276 = ~n_7273 &  n_7274;
assign n_7277 = ~n_7275 & ~n_7276;
assign n_7278 = ~x_2225 & ~n_7277;
assign n_7279 =  x_2225 & ~n_7276;
assign n_7280 = ~n_7275 &  n_7279;
assign n_7281 =  n_6534 & ~n_7280;
assign n_7282 = ~n_7278 &  n_7281;
assign n_7283 =  x_1393 &  n_6536;
assign n_7284 = ~x_2129 &  n_7254;
assign n_7285 =  x_2129 & ~n_7254;
assign n_7286 = ~n_7284 & ~n_7285;
assign n_7287 = ~n_7258 & ~n_7262;
assign n_7288 =  n_7286 & ~n_7287;
assign n_7289 = ~n_7286 &  n_7287;
assign n_7290 = ~n_7288 & ~n_7289;
assign n_7291 = ~x_561 & ~n_7290;
assign n_7292 =  x_561 & ~n_7289;
assign n_7293 = ~n_7288 &  n_7292;
assign n_7294 =  n_6531 & ~n_7293;
assign n_7295 = ~n_7291 &  n_7294;
assign n_7296 = ~n_7283 & ~n_7295;
assign n_7297 = ~n_7282 &  n_7296;
assign n_7298 =  x_1393 & ~n_7297;
assign n_7299 = ~x_1393 &  n_7297;
assign n_7300 = ~n_7298 & ~n_7299;
assign n_7301 = ~x_2736 &  n_7271;
assign n_7302 =  x_2736 & ~n_7271;
assign n_7303 = ~n_7301 & ~n_7302;
assign n_7304 = ~n_7275 & ~n_7279;
assign n_7305 =  n_7303 & ~n_7304;
assign n_7306 = ~n_7303 &  n_7304;
assign n_7307 = ~n_7305 & ~n_7306;
assign n_7308 = ~x_2224 & ~n_7307;
assign n_7309 =  x_2224 & ~n_7306;
assign n_7310 = ~n_7305 &  n_7309;
assign n_7311 =  n_6534 & ~n_7310;
assign n_7312 = ~n_7308 &  n_7311;
assign n_7313 =  x_1392 &  n_6536;
assign n_7314 = ~x_2128 &  n_7284;
assign n_7315 =  x_2128 & ~n_7284;
assign n_7316 = ~n_7314 & ~n_7315;
assign n_7317 = ~n_7288 & ~n_7292;
assign n_7318 =  n_7316 & ~n_7317;
assign n_7319 = ~n_7316 &  n_7317;
assign n_7320 = ~n_7318 & ~n_7319;
assign n_7321 = ~x_560 & ~n_7320;
assign n_7322 =  x_560 & ~n_7319;
assign n_7323 = ~n_7318 &  n_7322;
assign n_7324 =  n_6531 & ~n_7323;
assign n_7325 = ~n_7321 &  n_7324;
assign n_7326 = ~n_7313 & ~n_7325;
assign n_7327 = ~n_7312 &  n_7326;
assign n_7328 =  x_1392 & ~n_7327;
assign n_7329 = ~x_1392 &  n_7327;
assign n_7330 = ~n_7328 & ~n_7329;
assign n_7331 = ~x_2735 &  n_7301;
assign n_7332 =  x_2735 & ~n_7301;
assign n_7333 = ~n_7331 & ~n_7332;
assign n_7334 = ~n_7305 & ~n_7309;
assign n_7335 =  n_7333 & ~n_7334;
assign n_7336 = ~n_7333 &  n_7334;
assign n_7337 = ~n_7335 & ~n_7336;
assign n_7338 = ~x_2223 & ~n_7337;
assign n_7339 =  x_2223 & ~n_7336;
assign n_7340 = ~n_7335 &  n_7339;
assign n_7341 =  n_6534 & ~n_7340;
assign n_7342 = ~n_7338 &  n_7341;
assign n_7343 =  x_1391 &  n_6536;
assign n_7344 = ~x_2127 &  n_7314;
assign n_7345 =  x_2127 & ~n_7314;
assign n_7346 = ~n_7344 & ~n_7345;
assign n_7347 = ~n_7318 & ~n_7322;
assign n_7348 =  n_7346 & ~n_7347;
assign n_7349 = ~n_7346 &  n_7347;
assign n_7350 = ~n_7348 & ~n_7349;
assign n_7351 = ~x_559 & ~n_7350;
assign n_7352 =  x_559 & ~n_7349;
assign n_7353 = ~n_7348 &  n_7352;
assign n_7354 =  n_6531 & ~n_7353;
assign n_7355 = ~n_7351 &  n_7354;
assign n_7356 = ~n_7343 & ~n_7355;
assign n_7357 = ~n_7342 &  n_7356;
assign n_7358 =  x_1391 & ~n_7357;
assign n_7359 = ~x_1391 &  n_7357;
assign n_7360 = ~n_7358 & ~n_7359;
assign n_7361 = ~x_2734 &  n_7331;
assign n_7362 =  x_2734 & ~n_7331;
assign n_7363 = ~n_7361 & ~n_7362;
assign n_7364 = ~n_7335 & ~n_7339;
assign n_7365 =  n_7363 & ~n_7364;
assign n_7366 = ~n_7363 &  n_7364;
assign n_7367 = ~n_7365 & ~n_7366;
assign n_7368 = ~x_2222 & ~n_7367;
assign n_7369 =  x_2222 & ~n_7366;
assign n_7370 = ~n_7365 &  n_7369;
assign n_7371 =  n_6534 & ~n_7370;
assign n_7372 = ~n_7368 &  n_7371;
assign n_7373 =  x_1390 &  n_6536;
assign n_7374 = ~x_2126 &  n_7344;
assign n_7375 =  x_2126 & ~n_7344;
assign n_7376 = ~n_7374 & ~n_7375;
assign n_7377 = ~n_7348 & ~n_7352;
assign n_7378 =  n_7376 & ~n_7377;
assign n_7379 = ~n_7376 &  n_7377;
assign n_7380 = ~n_7378 & ~n_7379;
assign n_7381 = ~x_558 & ~n_7380;
assign n_7382 =  x_558 & ~n_7379;
assign n_7383 = ~n_7378 &  n_7382;
assign n_7384 =  n_6531 & ~n_7383;
assign n_7385 = ~n_7381 &  n_7384;
assign n_7386 = ~n_7373 & ~n_7385;
assign n_7387 = ~n_7372 &  n_7386;
assign n_7388 =  x_1390 & ~n_7387;
assign n_7389 = ~x_1390 &  n_7387;
assign n_7390 = ~n_7388 & ~n_7389;
assign n_7391 = ~x_2733 &  n_7361;
assign n_7392 =  x_2733 & ~n_7361;
assign n_7393 = ~n_7391 & ~n_7392;
assign n_7394 = ~n_7365 & ~n_7369;
assign n_7395 =  n_7393 & ~n_7394;
assign n_7396 = ~n_7393 &  n_7394;
assign n_7397 = ~n_7395 & ~n_7396;
assign n_7398 = ~x_2221 & ~n_7397;
assign n_7399 =  x_2221 & ~n_7396;
assign n_7400 = ~n_7395 &  n_7399;
assign n_7401 =  n_6534 & ~n_7400;
assign n_7402 = ~n_7398 &  n_7401;
assign n_7403 =  x_1389 &  n_6536;
assign n_7404 = ~x_2125 &  n_7374;
assign n_7405 =  x_2125 & ~n_7374;
assign n_7406 = ~n_7404 & ~n_7405;
assign n_7407 = ~n_7378 & ~n_7382;
assign n_7408 =  n_7406 & ~n_7407;
assign n_7409 = ~n_7406 &  n_7407;
assign n_7410 = ~n_7408 & ~n_7409;
assign n_7411 = ~x_557 & ~n_7410;
assign n_7412 =  x_557 & ~n_7409;
assign n_7413 = ~n_7408 &  n_7412;
assign n_7414 =  n_6531 & ~n_7413;
assign n_7415 = ~n_7411 &  n_7414;
assign n_7416 = ~n_7403 & ~n_7415;
assign n_7417 = ~n_7402 &  n_7416;
assign n_7418 =  x_1389 & ~n_7417;
assign n_7419 = ~x_1389 &  n_7417;
assign n_7420 = ~n_7418 & ~n_7419;
assign n_7421 = ~x_2732 &  n_7391;
assign n_7422 =  x_2732 & ~n_7391;
assign n_7423 = ~n_7421 & ~n_7422;
assign n_7424 = ~n_7395 & ~n_7399;
assign n_7425 =  n_7423 & ~n_7424;
assign n_7426 = ~n_7423 &  n_7424;
assign n_7427 = ~n_7425 & ~n_7426;
assign n_7428 = ~x_2220 & ~n_7427;
assign n_7429 =  x_2220 & ~n_7426;
assign n_7430 = ~n_7425 &  n_7429;
assign n_7431 =  n_6534 & ~n_7430;
assign n_7432 = ~n_7428 &  n_7431;
assign n_7433 =  x_1388 &  n_6536;
assign n_7434 = ~x_2124 &  n_7404;
assign n_7435 =  x_2124 & ~n_7404;
assign n_7436 = ~n_7434 & ~n_7435;
assign n_7437 = ~n_7408 & ~n_7412;
assign n_7438 =  n_7436 & ~n_7437;
assign n_7439 = ~n_7436 &  n_7437;
assign n_7440 = ~n_7438 & ~n_7439;
assign n_7441 = ~x_556 & ~n_7440;
assign n_7442 =  x_556 & ~n_7439;
assign n_7443 = ~n_7438 &  n_7442;
assign n_7444 =  n_6531 & ~n_7443;
assign n_7445 = ~n_7441 &  n_7444;
assign n_7446 = ~n_7433 & ~n_7445;
assign n_7447 = ~n_7432 &  n_7446;
assign n_7448 =  x_1388 & ~n_7447;
assign n_7449 = ~x_1388 &  n_7447;
assign n_7450 = ~n_7448 & ~n_7449;
assign n_7451 = ~n_7425 & ~n_7429;
assign n_7452 =  x_2219 & ~x_2731;
assign n_7453 = ~x_2219 &  x_2731;
assign n_7454 = ~n_7452 & ~n_7453;
assign n_7455 =  n_7421 &  n_7454;
assign n_7456 = ~n_7421 & ~n_7454;
assign n_7457 = ~n_7455 & ~n_7456;
assign n_7458 =  n_7451 & ~n_7457;
assign n_7459 = ~n_7451 &  n_7457;
assign n_7460 =  n_6534 & ~n_7459;
assign n_7461 = ~n_7458 &  n_7460;
assign n_7462 =  x_1387 &  n_6536;
assign n_7463 = ~n_7438 & ~n_7442;
assign n_7464 =  x_555 & ~x_2123;
assign n_7465 = ~x_555 &  x_2123;
assign n_7466 = ~n_7464 & ~n_7465;
assign n_7467 =  n_7434 &  n_7466;
assign n_7468 = ~n_7434 & ~n_7466;
assign n_7469 = ~n_7467 & ~n_7468;
assign n_7470 =  n_7463 & ~n_7469;
assign n_7471 = ~n_7463 &  n_7469;
assign n_7472 =  n_6531 & ~n_7471;
assign n_7473 = ~n_7470 &  n_7472;
assign n_7474 = ~n_7462 & ~n_7473;
assign n_7475 = ~n_7461 &  n_7474;
assign n_7476 =  x_1387 & ~n_7475;
assign n_7477 = ~x_1387 &  n_7475;
assign n_7478 = ~n_7476 & ~n_7477;
assign n_7479 =  n_980 &  n_3081;
assign n_7480 =  x_1386 & ~n_7479;
assign n_7481 =  i_32 &  n_7479;
assign n_7482 = ~n_7480 & ~n_7481;
assign n_7483 =  x_1386 & ~n_7482;
assign n_7484 = ~x_1386 &  n_7482;
assign n_7485 = ~n_7483 & ~n_7484;
assign n_7486 =  x_1385 & ~n_7479;
assign n_7487 =  i_31 &  n_7479;
assign n_7488 = ~n_7486 & ~n_7487;
assign n_7489 =  x_1385 & ~n_7488;
assign n_7490 = ~x_1385 &  n_7488;
assign n_7491 = ~n_7489 & ~n_7490;
assign n_7492 =  x_1384 & ~n_7479;
assign n_7493 =  i_30 &  n_7479;
assign n_7494 = ~n_7492 & ~n_7493;
assign n_7495 =  x_1384 & ~n_7494;
assign n_7496 = ~x_1384 &  n_7494;
assign n_7497 = ~n_7495 & ~n_7496;
assign n_7498 =  x_1383 & ~n_7479;
assign n_7499 =  i_29 &  n_7479;
assign n_7500 = ~n_7498 & ~n_7499;
assign n_7501 =  x_1383 & ~n_7500;
assign n_7502 = ~x_1383 &  n_7500;
assign n_7503 = ~n_7501 & ~n_7502;
assign n_7504 =  x_1382 & ~n_7479;
assign n_7505 =  i_28 &  n_7479;
assign n_7506 = ~n_7504 & ~n_7505;
assign n_7507 =  x_1382 & ~n_7506;
assign n_7508 = ~x_1382 &  n_7506;
assign n_7509 = ~n_7507 & ~n_7508;
assign n_7510 =  x_1381 & ~n_7479;
assign n_7511 =  i_27 &  n_7479;
assign n_7512 = ~n_7510 & ~n_7511;
assign n_7513 =  x_1381 & ~n_7512;
assign n_7514 = ~x_1381 &  n_7512;
assign n_7515 = ~n_7513 & ~n_7514;
assign n_7516 =  x_1380 & ~n_7479;
assign n_7517 =  i_26 &  n_7479;
assign n_7518 = ~n_7516 & ~n_7517;
assign n_7519 =  x_1380 & ~n_7518;
assign n_7520 = ~x_1380 &  n_7518;
assign n_7521 = ~n_7519 & ~n_7520;
assign n_7522 =  x_1379 & ~n_7479;
assign n_7523 =  i_25 &  n_7479;
assign n_7524 = ~n_7522 & ~n_7523;
assign n_7525 =  x_1379 & ~n_7524;
assign n_7526 = ~x_1379 &  n_7524;
assign n_7527 = ~n_7525 & ~n_7526;
assign n_7528 =  x_1378 & ~n_7479;
assign n_7529 =  i_24 &  n_7479;
assign n_7530 = ~n_7528 & ~n_7529;
assign n_7531 =  x_1378 & ~n_7530;
assign n_7532 = ~x_1378 &  n_7530;
assign n_7533 = ~n_7531 & ~n_7532;
assign n_7534 =  x_1377 & ~n_7479;
assign n_7535 =  i_23 &  n_7479;
assign n_7536 = ~n_7534 & ~n_7535;
assign n_7537 =  x_1377 & ~n_7536;
assign n_7538 = ~x_1377 &  n_7536;
assign n_7539 = ~n_7537 & ~n_7538;
assign n_7540 =  x_1376 & ~n_7479;
assign n_7541 =  i_22 &  n_7479;
assign n_7542 = ~n_7540 & ~n_7541;
assign n_7543 =  x_1376 & ~n_7542;
assign n_7544 = ~x_1376 &  n_7542;
assign n_7545 = ~n_7543 & ~n_7544;
assign n_7546 =  x_1375 & ~n_7479;
assign n_7547 =  i_21 &  n_7479;
assign n_7548 = ~n_7546 & ~n_7547;
assign n_7549 =  x_1375 & ~n_7548;
assign n_7550 = ~x_1375 &  n_7548;
assign n_7551 = ~n_7549 & ~n_7550;
assign n_7552 =  x_1374 & ~n_7479;
assign n_7553 =  i_20 &  n_7479;
assign n_7554 = ~n_7552 & ~n_7553;
assign n_7555 =  x_1374 & ~n_7554;
assign n_7556 = ~x_1374 &  n_7554;
assign n_7557 = ~n_7555 & ~n_7556;
assign n_7558 =  x_1373 & ~n_7479;
assign n_7559 =  i_19 &  n_7479;
assign n_7560 = ~n_7558 & ~n_7559;
assign n_7561 =  x_1373 & ~n_7560;
assign n_7562 = ~x_1373 &  n_7560;
assign n_7563 = ~n_7561 & ~n_7562;
assign n_7564 =  x_1372 & ~n_7479;
assign n_7565 =  i_18 &  n_7479;
assign n_7566 = ~n_7564 & ~n_7565;
assign n_7567 =  x_1372 & ~n_7566;
assign n_7568 = ~x_1372 &  n_7566;
assign n_7569 = ~n_7567 & ~n_7568;
assign n_7570 =  x_1371 & ~n_7479;
assign n_7571 =  i_17 &  n_7479;
assign n_7572 = ~n_7570 & ~n_7571;
assign n_7573 =  x_1371 & ~n_7572;
assign n_7574 = ~x_1371 &  n_7572;
assign n_7575 = ~n_7573 & ~n_7574;
assign n_7576 =  x_1370 & ~n_7479;
assign n_7577 =  i_16 &  n_7479;
assign n_7578 = ~n_7576 & ~n_7577;
assign n_7579 =  x_1370 & ~n_7578;
assign n_7580 = ~x_1370 &  n_7578;
assign n_7581 = ~n_7579 & ~n_7580;
assign n_7582 =  x_1369 & ~n_7479;
assign n_7583 =  i_15 &  n_7479;
assign n_7584 = ~n_7582 & ~n_7583;
assign n_7585 =  x_1369 & ~n_7584;
assign n_7586 = ~x_1369 &  n_7584;
assign n_7587 = ~n_7585 & ~n_7586;
assign n_7588 =  x_1368 & ~n_7479;
assign n_7589 =  i_14 &  n_7479;
assign n_7590 = ~n_7588 & ~n_7589;
assign n_7591 =  x_1368 & ~n_7590;
assign n_7592 = ~x_1368 &  n_7590;
assign n_7593 = ~n_7591 & ~n_7592;
assign n_7594 =  x_1367 & ~n_7479;
assign n_7595 =  i_13 &  n_7479;
assign n_7596 = ~n_7594 & ~n_7595;
assign n_7597 =  x_1367 & ~n_7596;
assign n_7598 = ~x_1367 &  n_7596;
assign n_7599 = ~n_7597 & ~n_7598;
assign n_7600 =  x_1366 & ~n_7479;
assign n_7601 =  i_12 &  n_7479;
assign n_7602 = ~n_7600 & ~n_7601;
assign n_7603 =  x_1366 & ~n_7602;
assign n_7604 = ~x_1366 &  n_7602;
assign n_7605 = ~n_7603 & ~n_7604;
assign n_7606 =  x_1365 & ~n_7479;
assign n_7607 =  i_11 &  n_7479;
assign n_7608 = ~n_7606 & ~n_7607;
assign n_7609 =  x_1365 & ~n_7608;
assign n_7610 = ~x_1365 &  n_7608;
assign n_7611 = ~n_7609 & ~n_7610;
assign n_7612 =  x_1364 & ~n_7479;
assign n_7613 =  i_10 &  n_7479;
assign n_7614 = ~n_7612 & ~n_7613;
assign n_7615 =  x_1364 & ~n_7614;
assign n_7616 = ~x_1364 &  n_7614;
assign n_7617 = ~n_7615 & ~n_7616;
assign n_7618 =  x_1363 & ~n_7479;
assign n_7619 =  i_9 &  n_7479;
assign n_7620 = ~n_7618 & ~n_7619;
assign n_7621 =  x_1363 & ~n_7620;
assign n_7622 = ~x_1363 &  n_7620;
assign n_7623 = ~n_7621 & ~n_7622;
assign n_7624 =  x_1362 & ~n_7479;
assign n_7625 =  i_8 &  n_7479;
assign n_7626 = ~n_7624 & ~n_7625;
assign n_7627 =  x_1362 & ~n_7626;
assign n_7628 = ~x_1362 &  n_7626;
assign n_7629 = ~n_7627 & ~n_7628;
assign n_7630 =  x_1361 & ~n_7479;
assign n_7631 =  i_7 &  n_7479;
assign n_7632 = ~n_7630 & ~n_7631;
assign n_7633 =  x_1361 & ~n_7632;
assign n_7634 = ~x_1361 &  n_7632;
assign n_7635 = ~n_7633 & ~n_7634;
assign n_7636 =  x_1360 & ~n_7479;
assign n_7637 =  i_6 &  n_7479;
assign n_7638 = ~n_7636 & ~n_7637;
assign n_7639 =  x_1360 & ~n_7638;
assign n_7640 = ~x_1360 &  n_7638;
assign n_7641 = ~n_7639 & ~n_7640;
assign n_7642 =  x_1359 & ~n_7479;
assign n_7643 =  i_5 &  n_7479;
assign n_7644 = ~n_7642 & ~n_7643;
assign n_7645 =  x_1359 & ~n_7644;
assign n_7646 = ~x_1359 &  n_7644;
assign n_7647 = ~n_7645 & ~n_7646;
assign n_7648 =  x_1358 & ~n_7479;
assign n_7649 =  i_4 &  n_7479;
assign n_7650 = ~n_7648 & ~n_7649;
assign n_7651 =  x_1358 & ~n_7650;
assign n_7652 = ~x_1358 &  n_7650;
assign n_7653 = ~n_7651 & ~n_7652;
assign n_7654 =  x_1357 & ~n_7479;
assign n_7655 =  i_3 &  n_7479;
assign n_7656 = ~n_7654 & ~n_7655;
assign n_7657 =  x_1357 & ~n_7656;
assign n_7658 = ~x_1357 &  n_7656;
assign n_7659 = ~n_7657 & ~n_7658;
assign n_7660 =  x_1356 & ~n_7479;
assign n_7661 =  i_2 &  n_7479;
assign n_7662 = ~n_7660 & ~n_7661;
assign n_7663 =  x_1356 & ~n_7662;
assign n_7664 = ~x_1356 &  n_7662;
assign n_7665 = ~n_7663 & ~n_7664;
assign n_7666 =  x_1355 & ~n_7479;
assign n_7667 =  i_1 &  n_7479;
assign n_7668 = ~n_7666 & ~n_7667;
assign n_7669 =  x_1355 & ~n_7668;
assign n_7670 = ~x_1355 &  n_7668;
assign n_7671 = ~n_7669 & ~n_7670;
assign n_7672 =  n_1707 &  n_6135;
assign n_7673 =  x_1354 & ~n_7672;
assign n_7674 =  i_32 &  n_7672;
assign n_7675 = ~n_7673 & ~n_7674;
assign n_7676 =  x_1354 & ~n_7675;
assign n_7677 = ~x_1354 &  n_7675;
assign n_7678 = ~n_7676 & ~n_7677;
assign n_7679 =  x_1353 & ~n_7672;
assign n_7680 =  i_31 &  n_7672;
assign n_7681 = ~n_7679 & ~n_7680;
assign n_7682 =  x_1353 & ~n_7681;
assign n_7683 = ~x_1353 &  n_7681;
assign n_7684 = ~n_7682 & ~n_7683;
assign n_7685 =  x_1352 & ~n_7672;
assign n_7686 =  i_30 &  n_7672;
assign n_7687 = ~n_7685 & ~n_7686;
assign n_7688 =  x_1352 & ~n_7687;
assign n_7689 = ~x_1352 &  n_7687;
assign n_7690 = ~n_7688 & ~n_7689;
assign n_7691 =  x_1351 & ~n_7672;
assign n_7692 =  i_29 &  n_7672;
assign n_7693 = ~n_7691 & ~n_7692;
assign n_7694 =  x_1351 & ~n_7693;
assign n_7695 = ~x_1351 &  n_7693;
assign n_7696 = ~n_7694 & ~n_7695;
assign n_7697 =  x_1350 & ~n_7672;
assign n_7698 =  i_28 &  n_7672;
assign n_7699 = ~n_7697 & ~n_7698;
assign n_7700 =  x_1350 & ~n_7699;
assign n_7701 = ~x_1350 &  n_7699;
assign n_7702 = ~n_7700 & ~n_7701;
assign n_7703 =  x_1349 & ~n_7672;
assign n_7704 =  i_27 &  n_7672;
assign n_7705 = ~n_7703 & ~n_7704;
assign n_7706 =  x_1349 & ~n_7705;
assign n_7707 = ~x_1349 &  n_7705;
assign n_7708 = ~n_7706 & ~n_7707;
assign n_7709 =  x_1348 & ~n_7672;
assign n_7710 =  i_26 &  n_7672;
assign n_7711 = ~n_7709 & ~n_7710;
assign n_7712 =  x_1348 & ~n_7711;
assign n_7713 = ~x_1348 &  n_7711;
assign n_7714 = ~n_7712 & ~n_7713;
assign n_7715 =  x_1347 & ~n_7672;
assign n_7716 =  i_25 &  n_7672;
assign n_7717 = ~n_7715 & ~n_7716;
assign n_7718 =  x_1347 & ~n_7717;
assign n_7719 = ~x_1347 &  n_7717;
assign n_7720 = ~n_7718 & ~n_7719;
assign n_7721 =  x_1346 & ~n_7672;
assign n_7722 =  i_24 &  n_7672;
assign n_7723 = ~n_7721 & ~n_7722;
assign n_7724 =  x_1346 & ~n_7723;
assign n_7725 = ~x_1346 &  n_7723;
assign n_7726 = ~n_7724 & ~n_7725;
assign n_7727 =  x_1345 & ~n_7672;
assign n_7728 =  i_23 &  n_7672;
assign n_7729 = ~n_7727 & ~n_7728;
assign n_7730 =  x_1345 & ~n_7729;
assign n_7731 = ~x_1345 &  n_7729;
assign n_7732 = ~n_7730 & ~n_7731;
assign n_7733 =  x_1344 & ~n_7672;
assign n_7734 =  i_22 &  n_7672;
assign n_7735 = ~n_7733 & ~n_7734;
assign n_7736 =  x_1344 & ~n_7735;
assign n_7737 = ~x_1344 &  n_7735;
assign n_7738 = ~n_7736 & ~n_7737;
assign n_7739 =  x_1343 & ~n_7672;
assign n_7740 =  i_21 &  n_7672;
assign n_7741 = ~n_7739 & ~n_7740;
assign n_7742 =  x_1343 & ~n_7741;
assign n_7743 = ~x_1343 &  n_7741;
assign n_7744 = ~n_7742 & ~n_7743;
assign n_7745 =  x_1342 & ~n_7672;
assign n_7746 =  i_20 &  n_7672;
assign n_7747 = ~n_7745 & ~n_7746;
assign n_7748 =  x_1342 & ~n_7747;
assign n_7749 = ~x_1342 &  n_7747;
assign n_7750 = ~n_7748 & ~n_7749;
assign n_7751 =  x_1341 & ~n_7672;
assign n_7752 =  i_19 &  n_7672;
assign n_7753 = ~n_7751 & ~n_7752;
assign n_7754 =  x_1341 & ~n_7753;
assign n_7755 = ~x_1341 &  n_7753;
assign n_7756 = ~n_7754 & ~n_7755;
assign n_7757 =  x_1340 & ~n_7672;
assign n_7758 =  i_18 &  n_7672;
assign n_7759 = ~n_7757 & ~n_7758;
assign n_7760 =  x_1340 & ~n_7759;
assign n_7761 = ~x_1340 &  n_7759;
assign n_7762 = ~n_7760 & ~n_7761;
assign n_7763 =  x_1339 & ~n_7672;
assign n_7764 =  i_17 &  n_7672;
assign n_7765 = ~n_7763 & ~n_7764;
assign n_7766 =  x_1339 & ~n_7765;
assign n_7767 = ~x_1339 &  n_7765;
assign n_7768 = ~n_7766 & ~n_7767;
assign n_7769 =  x_1338 & ~n_7672;
assign n_7770 =  i_16 &  n_7672;
assign n_7771 = ~n_7769 & ~n_7770;
assign n_7772 =  x_1338 & ~n_7771;
assign n_7773 = ~x_1338 &  n_7771;
assign n_7774 = ~n_7772 & ~n_7773;
assign n_7775 =  x_1337 & ~n_7672;
assign n_7776 =  i_15 &  n_7672;
assign n_7777 = ~n_7775 & ~n_7776;
assign n_7778 =  x_1337 & ~n_7777;
assign n_7779 = ~x_1337 &  n_7777;
assign n_7780 = ~n_7778 & ~n_7779;
assign n_7781 =  x_1336 & ~n_7672;
assign n_7782 =  i_14 &  n_7672;
assign n_7783 = ~n_7781 & ~n_7782;
assign n_7784 =  x_1336 & ~n_7783;
assign n_7785 = ~x_1336 &  n_7783;
assign n_7786 = ~n_7784 & ~n_7785;
assign n_7787 =  x_1335 & ~n_7672;
assign n_7788 =  i_13 &  n_7672;
assign n_7789 = ~n_7787 & ~n_7788;
assign n_7790 =  x_1335 & ~n_7789;
assign n_7791 = ~x_1335 &  n_7789;
assign n_7792 = ~n_7790 & ~n_7791;
assign n_7793 =  x_1334 & ~n_7672;
assign n_7794 =  i_12 &  n_7672;
assign n_7795 = ~n_7793 & ~n_7794;
assign n_7796 =  x_1334 & ~n_7795;
assign n_7797 = ~x_1334 &  n_7795;
assign n_7798 = ~n_7796 & ~n_7797;
assign n_7799 =  x_1333 & ~n_7672;
assign n_7800 =  i_11 &  n_7672;
assign n_7801 = ~n_7799 & ~n_7800;
assign n_7802 =  x_1333 & ~n_7801;
assign n_7803 = ~x_1333 &  n_7801;
assign n_7804 = ~n_7802 & ~n_7803;
assign n_7805 =  x_1332 & ~n_7672;
assign n_7806 =  i_10 &  n_7672;
assign n_7807 = ~n_7805 & ~n_7806;
assign n_7808 =  x_1332 & ~n_7807;
assign n_7809 = ~x_1332 &  n_7807;
assign n_7810 = ~n_7808 & ~n_7809;
assign n_7811 =  x_1331 & ~n_7672;
assign n_7812 =  i_9 &  n_7672;
assign n_7813 = ~n_7811 & ~n_7812;
assign n_7814 =  x_1331 & ~n_7813;
assign n_7815 = ~x_1331 &  n_7813;
assign n_7816 = ~n_7814 & ~n_7815;
assign n_7817 =  x_1330 & ~n_7672;
assign n_7818 =  i_8 &  n_7672;
assign n_7819 = ~n_7817 & ~n_7818;
assign n_7820 =  x_1330 & ~n_7819;
assign n_7821 = ~x_1330 &  n_7819;
assign n_7822 = ~n_7820 & ~n_7821;
assign n_7823 =  x_1329 & ~n_7672;
assign n_7824 =  i_7 &  n_7672;
assign n_7825 = ~n_7823 & ~n_7824;
assign n_7826 =  x_1329 & ~n_7825;
assign n_7827 = ~x_1329 &  n_7825;
assign n_7828 = ~n_7826 & ~n_7827;
assign n_7829 =  x_1328 & ~n_7672;
assign n_7830 =  i_6 &  n_7672;
assign n_7831 = ~n_7829 & ~n_7830;
assign n_7832 =  x_1328 & ~n_7831;
assign n_7833 = ~x_1328 &  n_7831;
assign n_7834 = ~n_7832 & ~n_7833;
assign n_7835 =  x_1327 & ~n_7672;
assign n_7836 =  i_5 &  n_7672;
assign n_7837 = ~n_7835 & ~n_7836;
assign n_7838 =  x_1327 & ~n_7837;
assign n_7839 = ~x_1327 &  n_7837;
assign n_7840 = ~n_7838 & ~n_7839;
assign n_7841 =  x_1326 & ~n_7672;
assign n_7842 =  i_4 &  n_7672;
assign n_7843 = ~n_7841 & ~n_7842;
assign n_7844 =  x_1326 & ~n_7843;
assign n_7845 = ~x_1326 &  n_7843;
assign n_7846 = ~n_7844 & ~n_7845;
assign n_7847 =  x_1325 & ~n_7672;
assign n_7848 =  i_3 &  n_7672;
assign n_7849 = ~n_7847 & ~n_7848;
assign n_7850 =  x_1325 & ~n_7849;
assign n_7851 = ~x_1325 &  n_7849;
assign n_7852 = ~n_7850 & ~n_7851;
assign n_7853 =  x_1324 & ~n_7672;
assign n_7854 =  i_2 &  n_7672;
assign n_7855 = ~n_7853 & ~n_7854;
assign n_7856 =  x_1324 & ~n_7855;
assign n_7857 = ~x_1324 &  n_7855;
assign n_7858 = ~n_7856 & ~n_7857;
assign n_7859 =  x_1323 & ~n_7672;
assign n_7860 =  i_1 &  n_7672;
assign n_7861 = ~n_7859 & ~n_7860;
assign n_7862 =  x_1323 & ~n_7861;
assign n_7863 = ~x_1323 &  n_7861;
assign n_7864 = ~n_7862 & ~n_7863;
assign n_7865 =  n_187 &  n_1178;
assign n_7866 =  n_6533 &  n_7865;
assign n_7867 =  x_1322 & ~n_7866;
assign n_7868 =  i_32 &  n_7866;
assign n_7869 = ~n_7867 & ~n_7868;
assign n_7870 =  x_1322 & ~n_7869;
assign n_7871 = ~x_1322 &  n_7869;
assign n_7872 = ~n_7870 & ~n_7871;
assign n_7873 =  x_1321 & ~n_7866;
assign n_7874 =  i_31 &  n_7866;
assign n_7875 = ~n_7873 & ~n_7874;
assign n_7876 =  x_1321 & ~n_7875;
assign n_7877 = ~x_1321 &  n_7875;
assign n_7878 = ~n_7876 & ~n_7877;
assign n_7879 =  x_1320 & ~n_7866;
assign n_7880 =  i_30 &  n_7866;
assign n_7881 = ~n_7879 & ~n_7880;
assign n_7882 =  x_1320 & ~n_7881;
assign n_7883 = ~x_1320 &  n_7881;
assign n_7884 = ~n_7882 & ~n_7883;
assign n_7885 =  x_1319 & ~n_7866;
assign n_7886 =  i_29 &  n_7866;
assign n_7887 = ~n_7885 & ~n_7886;
assign n_7888 =  x_1319 & ~n_7887;
assign n_7889 = ~x_1319 &  n_7887;
assign n_7890 = ~n_7888 & ~n_7889;
assign n_7891 =  x_1318 & ~n_7866;
assign n_7892 =  i_28 &  n_7866;
assign n_7893 = ~n_7891 & ~n_7892;
assign n_7894 =  x_1318 & ~n_7893;
assign n_7895 = ~x_1318 &  n_7893;
assign n_7896 = ~n_7894 & ~n_7895;
assign n_7897 =  x_1317 & ~n_7866;
assign n_7898 =  i_27 &  n_7866;
assign n_7899 = ~n_7897 & ~n_7898;
assign n_7900 =  x_1317 & ~n_7899;
assign n_7901 = ~x_1317 &  n_7899;
assign n_7902 = ~n_7900 & ~n_7901;
assign n_7903 =  x_1316 & ~n_7866;
assign n_7904 =  i_26 &  n_7866;
assign n_7905 = ~n_7903 & ~n_7904;
assign n_7906 =  x_1316 & ~n_7905;
assign n_7907 = ~x_1316 &  n_7905;
assign n_7908 = ~n_7906 & ~n_7907;
assign n_7909 =  x_1315 & ~n_7866;
assign n_7910 =  i_25 &  n_7866;
assign n_7911 = ~n_7909 & ~n_7910;
assign n_7912 =  x_1315 & ~n_7911;
assign n_7913 = ~x_1315 &  n_7911;
assign n_7914 = ~n_7912 & ~n_7913;
assign n_7915 =  x_1314 & ~n_7866;
assign n_7916 =  i_24 &  n_7866;
assign n_7917 = ~n_7915 & ~n_7916;
assign n_7918 =  x_1314 & ~n_7917;
assign n_7919 = ~x_1314 &  n_7917;
assign n_7920 = ~n_7918 & ~n_7919;
assign n_7921 =  x_1313 & ~n_7866;
assign n_7922 =  i_23 &  n_7866;
assign n_7923 = ~n_7921 & ~n_7922;
assign n_7924 =  x_1313 & ~n_7923;
assign n_7925 = ~x_1313 &  n_7923;
assign n_7926 = ~n_7924 & ~n_7925;
assign n_7927 =  x_1312 & ~n_7866;
assign n_7928 =  i_22 &  n_7866;
assign n_7929 = ~n_7927 & ~n_7928;
assign n_7930 =  x_1312 & ~n_7929;
assign n_7931 = ~x_1312 &  n_7929;
assign n_7932 = ~n_7930 & ~n_7931;
assign n_7933 =  x_1311 & ~n_7866;
assign n_7934 =  i_21 &  n_7866;
assign n_7935 = ~n_7933 & ~n_7934;
assign n_7936 =  x_1311 & ~n_7935;
assign n_7937 = ~x_1311 &  n_7935;
assign n_7938 = ~n_7936 & ~n_7937;
assign n_7939 =  x_1310 & ~n_7866;
assign n_7940 =  i_20 &  n_7866;
assign n_7941 = ~n_7939 & ~n_7940;
assign n_7942 =  x_1310 & ~n_7941;
assign n_7943 = ~x_1310 &  n_7941;
assign n_7944 = ~n_7942 & ~n_7943;
assign n_7945 =  x_1309 & ~n_7866;
assign n_7946 =  i_19 &  n_7866;
assign n_7947 = ~n_7945 & ~n_7946;
assign n_7948 =  x_1309 & ~n_7947;
assign n_7949 = ~x_1309 &  n_7947;
assign n_7950 = ~n_7948 & ~n_7949;
assign n_7951 =  x_1308 & ~n_7866;
assign n_7952 =  i_18 &  n_7866;
assign n_7953 = ~n_7951 & ~n_7952;
assign n_7954 =  x_1308 & ~n_7953;
assign n_7955 = ~x_1308 &  n_7953;
assign n_7956 = ~n_7954 & ~n_7955;
assign n_7957 =  x_1307 & ~n_7866;
assign n_7958 =  i_17 &  n_7866;
assign n_7959 = ~n_7957 & ~n_7958;
assign n_7960 =  x_1307 & ~n_7959;
assign n_7961 = ~x_1307 &  n_7959;
assign n_7962 = ~n_7960 & ~n_7961;
assign n_7963 =  x_1306 & ~n_7866;
assign n_7964 =  i_16 &  n_7866;
assign n_7965 = ~n_7963 & ~n_7964;
assign n_7966 =  x_1306 & ~n_7965;
assign n_7967 = ~x_1306 &  n_7965;
assign n_7968 = ~n_7966 & ~n_7967;
assign n_7969 =  x_1305 & ~n_7866;
assign n_7970 =  i_15 &  n_7866;
assign n_7971 = ~n_7969 & ~n_7970;
assign n_7972 =  x_1305 & ~n_7971;
assign n_7973 = ~x_1305 &  n_7971;
assign n_7974 = ~n_7972 & ~n_7973;
assign n_7975 =  x_1304 & ~n_7866;
assign n_7976 =  i_14 &  n_7866;
assign n_7977 = ~n_7975 & ~n_7976;
assign n_7978 =  x_1304 & ~n_7977;
assign n_7979 = ~x_1304 &  n_7977;
assign n_7980 = ~n_7978 & ~n_7979;
assign n_7981 =  x_1303 & ~n_7866;
assign n_7982 =  i_13 &  n_7866;
assign n_7983 = ~n_7981 & ~n_7982;
assign n_7984 =  x_1303 & ~n_7983;
assign n_7985 = ~x_1303 &  n_7983;
assign n_7986 = ~n_7984 & ~n_7985;
assign n_7987 =  x_1302 & ~n_7866;
assign n_7988 =  i_12 &  n_7866;
assign n_7989 = ~n_7987 & ~n_7988;
assign n_7990 =  x_1302 & ~n_7989;
assign n_7991 = ~x_1302 &  n_7989;
assign n_7992 = ~n_7990 & ~n_7991;
assign n_7993 =  x_1301 & ~n_7866;
assign n_7994 =  i_11 &  n_7866;
assign n_7995 = ~n_7993 & ~n_7994;
assign n_7996 =  x_1301 & ~n_7995;
assign n_7997 = ~x_1301 &  n_7995;
assign n_7998 = ~n_7996 & ~n_7997;
assign n_7999 =  x_1300 & ~n_7866;
assign n_8000 =  i_10 &  n_7866;
assign n_8001 = ~n_7999 & ~n_8000;
assign n_8002 =  x_1300 & ~n_8001;
assign n_8003 = ~x_1300 &  n_8001;
assign n_8004 = ~n_8002 & ~n_8003;
assign n_8005 =  x_1299 & ~n_7866;
assign n_8006 =  i_9 &  n_7866;
assign n_8007 = ~n_8005 & ~n_8006;
assign n_8008 =  x_1299 & ~n_8007;
assign n_8009 = ~x_1299 &  n_8007;
assign n_8010 = ~n_8008 & ~n_8009;
assign n_8011 =  x_1298 & ~n_7866;
assign n_8012 =  i_8 &  n_7866;
assign n_8013 = ~n_8011 & ~n_8012;
assign n_8014 =  x_1298 & ~n_8013;
assign n_8015 = ~x_1298 &  n_8013;
assign n_8016 = ~n_8014 & ~n_8015;
assign n_8017 =  x_1297 & ~n_7866;
assign n_8018 =  i_7 &  n_7866;
assign n_8019 = ~n_8017 & ~n_8018;
assign n_8020 =  x_1297 & ~n_8019;
assign n_8021 = ~x_1297 &  n_8019;
assign n_8022 = ~n_8020 & ~n_8021;
assign n_8023 =  x_1296 & ~n_7866;
assign n_8024 =  i_6 &  n_7866;
assign n_8025 = ~n_8023 & ~n_8024;
assign n_8026 =  x_1296 & ~n_8025;
assign n_8027 = ~x_1296 &  n_8025;
assign n_8028 = ~n_8026 & ~n_8027;
assign n_8029 =  x_1295 & ~n_7866;
assign n_8030 =  i_5 &  n_7866;
assign n_8031 = ~n_8029 & ~n_8030;
assign n_8032 =  x_1295 & ~n_8031;
assign n_8033 = ~x_1295 &  n_8031;
assign n_8034 = ~n_8032 & ~n_8033;
assign n_8035 =  x_1294 & ~n_7866;
assign n_8036 =  i_4 &  n_7866;
assign n_8037 = ~n_8035 & ~n_8036;
assign n_8038 =  x_1294 & ~n_8037;
assign n_8039 = ~x_1294 &  n_8037;
assign n_8040 = ~n_8038 & ~n_8039;
assign n_8041 =  x_1293 & ~n_7866;
assign n_8042 =  i_3 &  n_7866;
assign n_8043 = ~n_8041 & ~n_8042;
assign n_8044 =  x_1293 & ~n_8043;
assign n_8045 = ~x_1293 &  n_8043;
assign n_8046 = ~n_8044 & ~n_8045;
assign n_8047 =  x_1292 & ~n_7866;
assign n_8048 =  i_2 &  n_7866;
assign n_8049 = ~n_8047 & ~n_8048;
assign n_8050 =  x_1292 & ~n_8049;
assign n_8051 = ~x_1292 &  n_8049;
assign n_8052 = ~n_8050 & ~n_8051;
assign n_8053 =  x_1291 & ~n_7866;
assign n_8054 =  i_1 &  n_7866;
assign n_8055 = ~n_8053 & ~n_8054;
assign n_8056 =  x_1291 & ~n_8055;
assign n_8057 = ~x_1291 &  n_8055;
assign n_8058 = ~n_8056 & ~n_8057;
assign n_8059 =  x_41 &  n_2298;
assign n_8060 =  x_42 &  n_8059;
assign n_8061 =  n_8060 &  n_4057;
assign n_8062 =  x_1290 & ~n_8061;
assign n_8063 =  i_32 &  n_8061;
assign n_8064 = ~n_8062 & ~n_8063;
assign n_8065 =  x_1290 & ~n_8064;
assign n_8066 = ~x_1290 &  n_8064;
assign n_8067 = ~n_8065 & ~n_8066;
assign n_8068 =  x_1289 & ~n_8061;
assign n_8069 =  i_31 &  n_8061;
assign n_8070 = ~n_8068 & ~n_8069;
assign n_8071 =  x_1289 & ~n_8070;
assign n_8072 = ~x_1289 &  n_8070;
assign n_8073 = ~n_8071 & ~n_8072;
assign n_8074 =  x_1288 & ~n_8061;
assign n_8075 =  i_30 &  n_8061;
assign n_8076 = ~n_8074 & ~n_8075;
assign n_8077 =  x_1288 & ~n_8076;
assign n_8078 = ~x_1288 &  n_8076;
assign n_8079 = ~n_8077 & ~n_8078;
assign n_8080 =  x_1287 & ~n_8061;
assign n_8081 =  i_29 &  n_8061;
assign n_8082 = ~n_8080 & ~n_8081;
assign n_8083 =  x_1287 & ~n_8082;
assign n_8084 = ~x_1287 &  n_8082;
assign n_8085 = ~n_8083 & ~n_8084;
assign n_8086 =  x_1286 & ~n_8061;
assign n_8087 =  i_28 &  n_8061;
assign n_8088 = ~n_8086 & ~n_8087;
assign n_8089 =  x_1286 & ~n_8088;
assign n_8090 = ~x_1286 &  n_8088;
assign n_8091 = ~n_8089 & ~n_8090;
assign n_8092 =  x_1285 & ~n_8061;
assign n_8093 =  i_27 &  n_8061;
assign n_8094 = ~n_8092 & ~n_8093;
assign n_8095 =  x_1285 & ~n_8094;
assign n_8096 = ~x_1285 &  n_8094;
assign n_8097 = ~n_8095 & ~n_8096;
assign n_8098 =  x_1284 & ~n_8061;
assign n_8099 =  i_26 &  n_8061;
assign n_8100 = ~n_8098 & ~n_8099;
assign n_8101 =  x_1284 & ~n_8100;
assign n_8102 = ~x_1284 &  n_8100;
assign n_8103 = ~n_8101 & ~n_8102;
assign n_8104 =  x_1283 & ~n_8061;
assign n_8105 =  i_25 &  n_8061;
assign n_8106 = ~n_8104 & ~n_8105;
assign n_8107 =  x_1283 & ~n_8106;
assign n_8108 = ~x_1283 &  n_8106;
assign n_8109 = ~n_8107 & ~n_8108;
assign n_8110 =  x_1282 & ~n_8061;
assign n_8111 =  i_24 &  n_8061;
assign n_8112 = ~n_8110 & ~n_8111;
assign n_8113 =  x_1282 & ~n_8112;
assign n_8114 = ~x_1282 &  n_8112;
assign n_8115 = ~n_8113 & ~n_8114;
assign n_8116 =  x_1281 & ~n_8061;
assign n_8117 =  i_23 &  n_8061;
assign n_8118 = ~n_8116 & ~n_8117;
assign n_8119 =  x_1281 & ~n_8118;
assign n_8120 = ~x_1281 &  n_8118;
assign n_8121 = ~n_8119 & ~n_8120;
assign n_8122 =  x_1280 & ~n_8061;
assign n_8123 =  i_22 &  n_8061;
assign n_8124 = ~n_8122 & ~n_8123;
assign n_8125 =  x_1280 & ~n_8124;
assign n_8126 = ~x_1280 &  n_8124;
assign n_8127 = ~n_8125 & ~n_8126;
assign n_8128 =  x_1279 & ~n_8061;
assign n_8129 =  i_21 &  n_8061;
assign n_8130 = ~n_8128 & ~n_8129;
assign n_8131 =  x_1279 & ~n_8130;
assign n_8132 = ~x_1279 &  n_8130;
assign n_8133 = ~n_8131 & ~n_8132;
assign n_8134 =  x_1278 & ~n_8061;
assign n_8135 =  i_20 &  n_8061;
assign n_8136 = ~n_8134 & ~n_8135;
assign n_8137 =  x_1278 & ~n_8136;
assign n_8138 = ~x_1278 &  n_8136;
assign n_8139 = ~n_8137 & ~n_8138;
assign n_8140 =  x_1277 & ~n_8061;
assign n_8141 =  i_19 &  n_8061;
assign n_8142 = ~n_8140 & ~n_8141;
assign n_8143 =  x_1277 & ~n_8142;
assign n_8144 = ~x_1277 &  n_8142;
assign n_8145 = ~n_8143 & ~n_8144;
assign n_8146 =  x_1276 & ~n_8061;
assign n_8147 =  i_18 &  n_8061;
assign n_8148 = ~n_8146 & ~n_8147;
assign n_8149 =  x_1276 & ~n_8148;
assign n_8150 = ~x_1276 &  n_8148;
assign n_8151 = ~n_8149 & ~n_8150;
assign n_8152 =  x_1275 & ~n_8061;
assign n_8153 =  i_17 &  n_8061;
assign n_8154 = ~n_8152 & ~n_8153;
assign n_8155 =  x_1275 & ~n_8154;
assign n_8156 = ~x_1275 &  n_8154;
assign n_8157 = ~n_8155 & ~n_8156;
assign n_8158 =  x_1274 & ~n_8061;
assign n_8159 =  i_16 &  n_8061;
assign n_8160 = ~n_8158 & ~n_8159;
assign n_8161 =  x_1274 & ~n_8160;
assign n_8162 = ~x_1274 &  n_8160;
assign n_8163 = ~n_8161 & ~n_8162;
assign n_8164 =  x_1273 & ~n_8061;
assign n_8165 =  i_15 &  n_8061;
assign n_8166 = ~n_8164 & ~n_8165;
assign n_8167 =  x_1273 & ~n_8166;
assign n_8168 = ~x_1273 &  n_8166;
assign n_8169 = ~n_8167 & ~n_8168;
assign n_8170 =  x_1272 & ~n_8061;
assign n_8171 =  i_14 &  n_8061;
assign n_8172 = ~n_8170 & ~n_8171;
assign n_8173 =  x_1272 & ~n_8172;
assign n_8174 = ~x_1272 &  n_8172;
assign n_8175 = ~n_8173 & ~n_8174;
assign n_8176 =  x_1271 & ~n_8061;
assign n_8177 =  i_13 &  n_8061;
assign n_8178 = ~n_8176 & ~n_8177;
assign n_8179 =  x_1271 & ~n_8178;
assign n_8180 = ~x_1271 &  n_8178;
assign n_8181 = ~n_8179 & ~n_8180;
assign n_8182 =  x_1270 & ~n_8061;
assign n_8183 =  i_12 &  n_8061;
assign n_8184 = ~n_8182 & ~n_8183;
assign n_8185 =  x_1270 & ~n_8184;
assign n_8186 = ~x_1270 &  n_8184;
assign n_8187 = ~n_8185 & ~n_8186;
assign n_8188 =  x_1269 & ~n_8061;
assign n_8189 =  i_11 &  n_8061;
assign n_8190 = ~n_8188 & ~n_8189;
assign n_8191 =  x_1269 & ~n_8190;
assign n_8192 = ~x_1269 &  n_8190;
assign n_8193 = ~n_8191 & ~n_8192;
assign n_8194 =  x_1268 & ~n_8061;
assign n_8195 =  i_10 &  n_8061;
assign n_8196 = ~n_8194 & ~n_8195;
assign n_8197 =  x_1268 & ~n_8196;
assign n_8198 = ~x_1268 &  n_8196;
assign n_8199 = ~n_8197 & ~n_8198;
assign n_8200 =  x_1267 & ~n_8061;
assign n_8201 =  i_9 &  n_8061;
assign n_8202 = ~n_8200 & ~n_8201;
assign n_8203 =  x_1267 & ~n_8202;
assign n_8204 = ~x_1267 &  n_8202;
assign n_8205 = ~n_8203 & ~n_8204;
assign n_8206 =  x_1266 & ~n_8061;
assign n_8207 =  i_8 &  n_8061;
assign n_8208 = ~n_8206 & ~n_8207;
assign n_8209 =  x_1266 & ~n_8208;
assign n_8210 = ~x_1266 &  n_8208;
assign n_8211 = ~n_8209 & ~n_8210;
assign n_8212 =  x_1265 & ~n_8061;
assign n_8213 =  i_7 &  n_8061;
assign n_8214 = ~n_8212 & ~n_8213;
assign n_8215 =  x_1265 & ~n_8214;
assign n_8216 = ~x_1265 &  n_8214;
assign n_8217 = ~n_8215 & ~n_8216;
assign n_8218 =  x_1264 & ~n_8061;
assign n_8219 =  i_6 &  n_8061;
assign n_8220 = ~n_8218 & ~n_8219;
assign n_8221 =  x_1264 & ~n_8220;
assign n_8222 = ~x_1264 &  n_8220;
assign n_8223 = ~n_8221 & ~n_8222;
assign n_8224 =  x_1263 & ~n_8061;
assign n_8225 =  i_5 &  n_8061;
assign n_8226 = ~n_8224 & ~n_8225;
assign n_8227 =  x_1263 & ~n_8226;
assign n_8228 = ~x_1263 &  n_8226;
assign n_8229 = ~n_8227 & ~n_8228;
assign n_8230 =  x_1262 & ~n_8061;
assign n_8231 =  i_4 &  n_8061;
assign n_8232 = ~n_8230 & ~n_8231;
assign n_8233 =  x_1262 & ~n_8232;
assign n_8234 = ~x_1262 &  n_8232;
assign n_8235 = ~n_8233 & ~n_8234;
assign n_8236 =  x_1261 & ~n_8061;
assign n_8237 =  i_3 &  n_8061;
assign n_8238 = ~n_8236 & ~n_8237;
assign n_8239 =  x_1261 & ~n_8238;
assign n_8240 = ~x_1261 &  n_8238;
assign n_8241 = ~n_8239 & ~n_8240;
assign n_8242 =  x_1260 & ~n_8061;
assign n_8243 =  i_2 &  n_8061;
assign n_8244 = ~n_8242 & ~n_8243;
assign n_8245 =  x_1260 & ~n_8244;
assign n_8246 = ~x_1260 &  n_8244;
assign n_8247 = ~n_8245 & ~n_8246;
assign n_8248 =  x_1259 & ~n_8061;
assign n_8249 =  i_1 &  n_8061;
assign n_8250 = ~n_8248 & ~n_8249;
assign n_8251 =  x_1259 & ~n_8250;
assign n_8252 = ~x_1259 &  n_8250;
assign n_8253 = ~n_8251 & ~n_8252;
assign n_8254 =  n_1706 &  n_2298;
assign n_8255 =  n_389 &  n_8254;
assign n_8256 =  n_190 &  n_8255;
assign n_8257 =  x_1258 & ~n_8256;
assign n_8258 =  i_32 &  n_8256;
assign n_8259 = ~n_8257 & ~n_8258;
assign n_8260 =  x_1258 & ~n_8259;
assign n_8261 = ~x_1258 &  n_8259;
assign n_8262 = ~n_8260 & ~n_8261;
assign n_8263 =  x_1257 & ~n_8256;
assign n_8264 =  i_31 &  n_8256;
assign n_8265 = ~n_8263 & ~n_8264;
assign n_8266 =  x_1257 & ~n_8265;
assign n_8267 = ~x_1257 &  n_8265;
assign n_8268 = ~n_8266 & ~n_8267;
assign n_8269 =  x_1256 & ~n_8256;
assign n_8270 =  i_30 &  n_8256;
assign n_8271 = ~n_8269 & ~n_8270;
assign n_8272 =  x_1256 & ~n_8271;
assign n_8273 = ~x_1256 &  n_8271;
assign n_8274 = ~n_8272 & ~n_8273;
assign n_8275 =  x_1255 & ~n_8256;
assign n_8276 =  i_29 &  n_8256;
assign n_8277 = ~n_8275 & ~n_8276;
assign n_8278 =  x_1255 & ~n_8277;
assign n_8279 = ~x_1255 &  n_8277;
assign n_8280 = ~n_8278 & ~n_8279;
assign n_8281 =  x_1254 & ~n_8256;
assign n_8282 =  i_28 &  n_8256;
assign n_8283 = ~n_8281 & ~n_8282;
assign n_8284 =  x_1254 & ~n_8283;
assign n_8285 = ~x_1254 &  n_8283;
assign n_8286 = ~n_8284 & ~n_8285;
assign n_8287 =  x_1253 & ~n_8256;
assign n_8288 =  i_27 &  n_8256;
assign n_8289 = ~n_8287 & ~n_8288;
assign n_8290 =  x_1253 & ~n_8289;
assign n_8291 = ~x_1253 &  n_8289;
assign n_8292 = ~n_8290 & ~n_8291;
assign n_8293 =  x_1252 & ~n_8256;
assign n_8294 =  i_26 &  n_8256;
assign n_8295 = ~n_8293 & ~n_8294;
assign n_8296 =  x_1252 & ~n_8295;
assign n_8297 = ~x_1252 &  n_8295;
assign n_8298 = ~n_8296 & ~n_8297;
assign n_8299 =  x_1251 & ~n_8256;
assign n_8300 =  i_25 &  n_8256;
assign n_8301 = ~n_8299 & ~n_8300;
assign n_8302 =  x_1251 & ~n_8301;
assign n_8303 = ~x_1251 &  n_8301;
assign n_8304 = ~n_8302 & ~n_8303;
assign n_8305 =  x_1250 & ~n_8256;
assign n_8306 =  i_24 &  n_8256;
assign n_8307 = ~n_8305 & ~n_8306;
assign n_8308 =  x_1250 & ~n_8307;
assign n_8309 = ~x_1250 &  n_8307;
assign n_8310 = ~n_8308 & ~n_8309;
assign n_8311 =  x_1249 & ~n_8256;
assign n_8312 =  i_23 &  n_8256;
assign n_8313 = ~n_8311 & ~n_8312;
assign n_8314 =  x_1249 & ~n_8313;
assign n_8315 = ~x_1249 &  n_8313;
assign n_8316 = ~n_8314 & ~n_8315;
assign n_8317 =  x_1248 & ~n_8256;
assign n_8318 =  i_22 &  n_8256;
assign n_8319 = ~n_8317 & ~n_8318;
assign n_8320 =  x_1248 & ~n_8319;
assign n_8321 = ~x_1248 &  n_8319;
assign n_8322 = ~n_8320 & ~n_8321;
assign n_8323 =  x_1247 & ~n_8256;
assign n_8324 =  i_21 &  n_8256;
assign n_8325 = ~n_8323 & ~n_8324;
assign n_8326 =  x_1247 & ~n_8325;
assign n_8327 = ~x_1247 &  n_8325;
assign n_8328 = ~n_8326 & ~n_8327;
assign n_8329 =  x_1246 & ~n_8256;
assign n_8330 =  i_20 &  n_8256;
assign n_8331 = ~n_8329 & ~n_8330;
assign n_8332 =  x_1246 & ~n_8331;
assign n_8333 = ~x_1246 &  n_8331;
assign n_8334 = ~n_8332 & ~n_8333;
assign n_8335 =  x_1245 & ~n_8256;
assign n_8336 =  i_19 &  n_8256;
assign n_8337 = ~n_8335 & ~n_8336;
assign n_8338 =  x_1245 & ~n_8337;
assign n_8339 = ~x_1245 &  n_8337;
assign n_8340 = ~n_8338 & ~n_8339;
assign n_8341 =  x_1244 & ~n_8256;
assign n_8342 =  i_18 &  n_8256;
assign n_8343 = ~n_8341 & ~n_8342;
assign n_8344 =  x_1244 & ~n_8343;
assign n_8345 = ~x_1244 &  n_8343;
assign n_8346 = ~n_8344 & ~n_8345;
assign n_8347 =  x_1243 & ~n_8256;
assign n_8348 =  i_17 &  n_8256;
assign n_8349 = ~n_8347 & ~n_8348;
assign n_8350 =  x_1243 & ~n_8349;
assign n_8351 = ~x_1243 &  n_8349;
assign n_8352 = ~n_8350 & ~n_8351;
assign n_8353 =  x_1242 & ~n_8256;
assign n_8354 =  i_16 &  n_8256;
assign n_8355 = ~n_8353 & ~n_8354;
assign n_8356 =  x_1242 & ~n_8355;
assign n_8357 = ~x_1242 &  n_8355;
assign n_8358 = ~n_8356 & ~n_8357;
assign n_8359 =  x_1241 & ~n_8256;
assign n_8360 =  i_15 &  n_8256;
assign n_8361 = ~n_8359 & ~n_8360;
assign n_8362 =  x_1241 & ~n_8361;
assign n_8363 = ~x_1241 &  n_8361;
assign n_8364 = ~n_8362 & ~n_8363;
assign n_8365 =  x_1240 & ~n_8256;
assign n_8366 =  i_14 &  n_8256;
assign n_8367 = ~n_8365 & ~n_8366;
assign n_8368 =  x_1240 & ~n_8367;
assign n_8369 = ~x_1240 &  n_8367;
assign n_8370 = ~n_8368 & ~n_8369;
assign n_8371 =  x_1239 & ~n_8256;
assign n_8372 =  i_13 &  n_8256;
assign n_8373 = ~n_8371 & ~n_8372;
assign n_8374 =  x_1239 & ~n_8373;
assign n_8375 = ~x_1239 &  n_8373;
assign n_8376 = ~n_8374 & ~n_8375;
assign n_8377 =  x_1238 & ~n_8256;
assign n_8378 =  i_12 &  n_8256;
assign n_8379 = ~n_8377 & ~n_8378;
assign n_8380 =  x_1238 & ~n_8379;
assign n_8381 = ~x_1238 &  n_8379;
assign n_8382 = ~n_8380 & ~n_8381;
assign n_8383 =  x_1237 & ~n_8256;
assign n_8384 =  i_11 &  n_8256;
assign n_8385 = ~n_8383 & ~n_8384;
assign n_8386 =  x_1237 & ~n_8385;
assign n_8387 = ~x_1237 &  n_8385;
assign n_8388 = ~n_8386 & ~n_8387;
assign n_8389 =  x_1236 & ~n_8256;
assign n_8390 =  i_10 &  n_8256;
assign n_8391 = ~n_8389 & ~n_8390;
assign n_8392 =  x_1236 & ~n_8391;
assign n_8393 = ~x_1236 &  n_8391;
assign n_8394 = ~n_8392 & ~n_8393;
assign n_8395 =  x_1235 & ~n_8256;
assign n_8396 =  i_9 &  n_8256;
assign n_8397 = ~n_8395 & ~n_8396;
assign n_8398 =  x_1235 & ~n_8397;
assign n_8399 = ~x_1235 &  n_8397;
assign n_8400 = ~n_8398 & ~n_8399;
assign n_8401 =  x_1234 & ~n_8256;
assign n_8402 =  i_8 &  n_8256;
assign n_8403 = ~n_8401 & ~n_8402;
assign n_8404 =  x_1234 & ~n_8403;
assign n_8405 = ~x_1234 &  n_8403;
assign n_8406 = ~n_8404 & ~n_8405;
assign n_8407 =  x_1233 & ~n_8256;
assign n_8408 =  i_7 &  n_8256;
assign n_8409 = ~n_8407 & ~n_8408;
assign n_8410 =  x_1233 & ~n_8409;
assign n_8411 = ~x_1233 &  n_8409;
assign n_8412 = ~n_8410 & ~n_8411;
assign n_8413 =  x_1232 & ~n_8256;
assign n_8414 =  i_6 &  n_8256;
assign n_8415 = ~n_8413 & ~n_8414;
assign n_8416 =  x_1232 & ~n_8415;
assign n_8417 = ~x_1232 &  n_8415;
assign n_8418 = ~n_8416 & ~n_8417;
assign n_8419 =  x_1231 & ~n_8256;
assign n_8420 =  i_5 &  n_8256;
assign n_8421 = ~n_8419 & ~n_8420;
assign n_8422 =  x_1231 & ~n_8421;
assign n_8423 = ~x_1231 &  n_8421;
assign n_8424 = ~n_8422 & ~n_8423;
assign n_8425 =  x_1230 & ~n_8256;
assign n_8426 =  i_4 &  n_8256;
assign n_8427 = ~n_8425 & ~n_8426;
assign n_8428 =  x_1230 & ~n_8427;
assign n_8429 = ~x_1230 &  n_8427;
assign n_8430 = ~n_8428 & ~n_8429;
assign n_8431 =  x_1229 & ~n_8256;
assign n_8432 =  i_3 &  n_8256;
assign n_8433 = ~n_8431 & ~n_8432;
assign n_8434 =  x_1229 & ~n_8433;
assign n_8435 = ~x_1229 &  n_8433;
assign n_8436 = ~n_8434 & ~n_8435;
assign n_8437 =  x_1228 & ~n_8256;
assign n_8438 =  i_2 &  n_8256;
assign n_8439 = ~n_8437 & ~n_8438;
assign n_8440 =  x_1228 & ~n_8439;
assign n_8441 = ~x_1228 &  n_8439;
assign n_8442 = ~n_8440 & ~n_8441;
assign n_8443 =  x_1227 & ~n_8256;
assign n_8444 =  i_1 &  n_8256;
assign n_8445 = ~n_8443 & ~n_8444;
assign n_8446 =  x_1227 & ~n_8445;
assign n_8447 = ~x_1227 &  n_8445;
assign n_8448 = ~n_8446 & ~n_8447;
assign n_8449 =  n_1707 &  n_390;
assign n_8450 =  x_1226 & ~n_8449;
assign n_8451 =  i_32 &  n_8449;
assign n_8452 = ~n_8450 & ~n_8451;
assign n_8453 =  x_1226 & ~n_8452;
assign n_8454 = ~x_1226 &  n_8452;
assign n_8455 = ~n_8453 & ~n_8454;
assign n_8456 =  x_1225 & ~n_8449;
assign n_8457 =  i_31 &  n_8449;
assign n_8458 = ~n_8456 & ~n_8457;
assign n_8459 =  x_1225 & ~n_8458;
assign n_8460 = ~x_1225 &  n_8458;
assign n_8461 = ~n_8459 & ~n_8460;
assign n_8462 =  x_1224 & ~n_8449;
assign n_8463 =  i_30 &  n_8449;
assign n_8464 = ~n_8462 & ~n_8463;
assign n_8465 =  x_1224 & ~n_8464;
assign n_8466 = ~x_1224 &  n_8464;
assign n_8467 = ~n_8465 & ~n_8466;
assign n_8468 =  x_1223 & ~n_8449;
assign n_8469 =  i_29 &  n_8449;
assign n_8470 = ~n_8468 & ~n_8469;
assign n_8471 =  x_1223 & ~n_8470;
assign n_8472 = ~x_1223 &  n_8470;
assign n_8473 = ~n_8471 & ~n_8472;
assign n_8474 =  x_1222 & ~n_8449;
assign n_8475 =  i_28 &  n_8449;
assign n_8476 = ~n_8474 & ~n_8475;
assign n_8477 =  x_1222 & ~n_8476;
assign n_8478 = ~x_1222 &  n_8476;
assign n_8479 = ~n_8477 & ~n_8478;
assign n_8480 =  x_1221 & ~n_8449;
assign n_8481 =  i_27 &  n_8449;
assign n_8482 = ~n_8480 & ~n_8481;
assign n_8483 =  x_1221 & ~n_8482;
assign n_8484 = ~x_1221 &  n_8482;
assign n_8485 = ~n_8483 & ~n_8484;
assign n_8486 =  x_1220 & ~n_8449;
assign n_8487 =  i_26 &  n_8449;
assign n_8488 = ~n_8486 & ~n_8487;
assign n_8489 =  x_1220 & ~n_8488;
assign n_8490 = ~x_1220 &  n_8488;
assign n_8491 = ~n_8489 & ~n_8490;
assign n_8492 =  x_1219 & ~n_8449;
assign n_8493 =  i_25 &  n_8449;
assign n_8494 = ~n_8492 & ~n_8493;
assign n_8495 =  x_1219 & ~n_8494;
assign n_8496 = ~x_1219 &  n_8494;
assign n_8497 = ~n_8495 & ~n_8496;
assign n_8498 =  x_1218 & ~n_8449;
assign n_8499 =  i_24 &  n_8449;
assign n_8500 = ~n_8498 & ~n_8499;
assign n_8501 =  x_1218 & ~n_8500;
assign n_8502 = ~x_1218 &  n_8500;
assign n_8503 = ~n_8501 & ~n_8502;
assign n_8504 =  x_1217 & ~n_8449;
assign n_8505 =  i_23 &  n_8449;
assign n_8506 = ~n_8504 & ~n_8505;
assign n_8507 =  x_1217 & ~n_8506;
assign n_8508 = ~x_1217 &  n_8506;
assign n_8509 = ~n_8507 & ~n_8508;
assign n_8510 =  x_1216 & ~n_8449;
assign n_8511 =  i_22 &  n_8449;
assign n_8512 = ~n_8510 & ~n_8511;
assign n_8513 =  x_1216 & ~n_8512;
assign n_8514 = ~x_1216 &  n_8512;
assign n_8515 = ~n_8513 & ~n_8514;
assign n_8516 =  x_1215 & ~n_8449;
assign n_8517 =  i_21 &  n_8449;
assign n_8518 = ~n_8516 & ~n_8517;
assign n_8519 =  x_1215 & ~n_8518;
assign n_8520 = ~x_1215 &  n_8518;
assign n_8521 = ~n_8519 & ~n_8520;
assign n_8522 =  x_1214 & ~n_8449;
assign n_8523 =  i_20 &  n_8449;
assign n_8524 = ~n_8522 & ~n_8523;
assign n_8525 =  x_1214 & ~n_8524;
assign n_8526 = ~x_1214 &  n_8524;
assign n_8527 = ~n_8525 & ~n_8526;
assign n_8528 =  x_1213 & ~n_8449;
assign n_8529 =  i_19 &  n_8449;
assign n_8530 = ~n_8528 & ~n_8529;
assign n_8531 =  x_1213 & ~n_8530;
assign n_8532 = ~x_1213 &  n_8530;
assign n_8533 = ~n_8531 & ~n_8532;
assign n_8534 =  x_1212 & ~n_8449;
assign n_8535 =  i_18 &  n_8449;
assign n_8536 = ~n_8534 & ~n_8535;
assign n_8537 =  x_1212 & ~n_8536;
assign n_8538 = ~x_1212 &  n_8536;
assign n_8539 = ~n_8537 & ~n_8538;
assign n_8540 =  x_1211 & ~n_8449;
assign n_8541 =  i_17 &  n_8449;
assign n_8542 = ~n_8540 & ~n_8541;
assign n_8543 =  x_1211 & ~n_8542;
assign n_8544 = ~x_1211 &  n_8542;
assign n_8545 = ~n_8543 & ~n_8544;
assign n_8546 =  x_1210 & ~n_8449;
assign n_8547 =  i_16 &  n_8449;
assign n_8548 = ~n_8546 & ~n_8547;
assign n_8549 =  x_1210 & ~n_8548;
assign n_8550 = ~x_1210 &  n_8548;
assign n_8551 = ~n_8549 & ~n_8550;
assign n_8552 =  x_1209 & ~n_8449;
assign n_8553 =  i_15 &  n_8449;
assign n_8554 = ~n_8552 & ~n_8553;
assign n_8555 =  x_1209 & ~n_8554;
assign n_8556 = ~x_1209 &  n_8554;
assign n_8557 = ~n_8555 & ~n_8556;
assign n_8558 =  x_1208 & ~n_8449;
assign n_8559 =  i_14 &  n_8449;
assign n_8560 = ~n_8558 & ~n_8559;
assign n_8561 =  x_1208 & ~n_8560;
assign n_8562 = ~x_1208 &  n_8560;
assign n_8563 = ~n_8561 & ~n_8562;
assign n_8564 =  x_1207 & ~n_8449;
assign n_8565 =  i_13 &  n_8449;
assign n_8566 = ~n_8564 & ~n_8565;
assign n_8567 =  x_1207 & ~n_8566;
assign n_8568 = ~x_1207 &  n_8566;
assign n_8569 = ~n_8567 & ~n_8568;
assign n_8570 =  x_1206 & ~n_8449;
assign n_8571 =  i_12 &  n_8449;
assign n_8572 = ~n_8570 & ~n_8571;
assign n_8573 =  x_1206 & ~n_8572;
assign n_8574 = ~x_1206 &  n_8572;
assign n_8575 = ~n_8573 & ~n_8574;
assign n_8576 =  x_1205 & ~n_8449;
assign n_8577 =  i_11 &  n_8449;
assign n_8578 = ~n_8576 & ~n_8577;
assign n_8579 =  x_1205 & ~n_8578;
assign n_8580 = ~x_1205 &  n_8578;
assign n_8581 = ~n_8579 & ~n_8580;
assign n_8582 =  x_1204 & ~n_8449;
assign n_8583 =  i_10 &  n_8449;
assign n_8584 = ~n_8582 & ~n_8583;
assign n_8585 =  x_1204 & ~n_8584;
assign n_8586 = ~x_1204 &  n_8584;
assign n_8587 = ~n_8585 & ~n_8586;
assign n_8588 =  x_1203 & ~n_8449;
assign n_8589 =  i_9 &  n_8449;
assign n_8590 = ~n_8588 & ~n_8589;
assign n_8591 =  x_1203 & ~n_8590;
assign n_8592 = ~x_1203 &  n_8590;
assign n_8593 = ~n_8591 & ~n_8592;
assign n_8594 =  x_1202 & ~n_8449;
assign n_8595 =  i_8 &  n_8449;
assign n_8596 = ~n_8594 & ~n_8595;
assign n_8597 =  x_1202 & ~n_8596;
assign n_8598 = ~x_1202 &  n_8596;
assign n_8599 = ~n_8597 & ~n_8598;
assign n_8600 =  x_1201 & ~n_8449;
assign n_8601 =  i_7 &  n_8449;
assign n_8602 = ~n_8600 & ~n_8601;
assign n_8603 =  x_1201 & ~n_8602;
assign n_8604 = ~x_1201 &  n_8602;
assign n_8605 = ~n_8603 & ~n_8604;
assign n_8606 =  x_1200 & ~n_8449;
assign n_8607 =  i_6 &  n_8449;
assign n_8608 = ~n_8606 & ~n_8607;
assign n_8609 =  x_1200 & ~n_8608;
assign n_8610 = ~x_1200 &  n_8608;
assign n_8611 = ~n_8609 & ~n_8610;
assign n_8612 =  x_1199 & ~n_8449;
assign n_8613 =  i_5 &  n_8449;
assign n_8614 = ~n_8612 & ~n_8613;
assign n_8615 =  x_1199 & ~n_8614;
assign n_8616 = ~x_1199 &  n_8614;
assign n_8617 = ~n_8615 & ~n_8616;
assign n_8618 =  x_1198 & ~n_8449;
assign n_8619 =  i_4 &  n_8449;
assign n_8620 = ~n_8618 & ~n_8619;
assign n_8621 =  x_1198 & ~n_8620;
assign n_8622 = ~x_1198 &  n_8620;
assign n_8623 = ~n_8621 & ~n_8622;
assign n_8624 =  x_1197 & ~n_8449;
assign n_8625 =  i_3 &  n_8449;
assign n_8626 = ~n_8624 & ~n_8625;
assign n_8627 =  x_1197 & ~n_8626;
assign n_8628 = ~x_1197 &  n_8626;
assign n_8629 = ~n_8627 & ~n_8628;
assign n_8630 =  x_1196 & ~n_8449;
assign n_8631 =  i_2 &  n_8449;
assign n_8632 = ~n_8630 & ~n_8631;
assign n_8633 =  x_1196 & ~n_8632;
assign n_8634 = ~x_1196 &  n_8632;
assign n_8635 = ~n_8633 & ~n_8634;
assign n_8636 =  x_1195 & ~n_8449;
assign n_8637 =  i_1 &  n_8449;
assign n_8638 = ~n_8636 & ~n_8637;
assign n_8639 =  x_1195 & ~n_8638;
assign n_8640 = ~x_1195 &  n_8638;
assign n_8641 = ~n_8639 & ~n_8640;
assign n_8642 =  x_1194 & ~n_984;
assign n_8643 = ~n_985 & ~n_8642;
assign n_8644 =  x_1194 & ~n_8643;
assign n_8645 = ~x_1194 &  n_8643;
assign n_8646 = ~n_8644 & ~n_8645;
assign n_8647 =  x_1193 & ~n_984;
assign n_8648 = ~n_991 & ~n_8647;
assign n_8649 =  x_1193 & ~n_8648;
assign n_8650 = ~x_1193 &  n_8648;
assign n_8651 = ~n_8649 & ~n_8650;
assign n_8652 =  x_1192 & ~n_984;
assign n_8653 = ~n_997 & ~n_8652;
assign n_8654 =  x_1192 & ~n_8653;
assign n_8655 = ~x_1192 &  n_8653;
assign n_8656 = ~n_8654 & ~n_8655;
assign n_8657 =  x_1191 & ~n_984;
assign n_8658 = ~n_1003 & ~n_8657;
assign n_8659 =  x_1191 & ~n_8658;
assign n_8660 = ~x_1191 &  n_8658;
assign n_8661 = ~n_8659 & ~n_8660;
assign n_8662 =  x_1190 & ~n_984;
assign n_8663 = ~n_1009 & ~n_8662;
assign n_8664 =  x_1190 & ~n_8663;
assign n_8665 = ~x_1190 &  n_8663;
assign n_8666 = ~n_8664 & ~n_8665;
assign n_8667 =  x_1189 & ~n_984;
assign n_8668 = ~n_1015 & ~n_8667;
assign n_8669 =  x_1189 & ~n_8668;
assign n_8670 = ~x_1189 &  n_8668;
assign n_8671 = ~n_8669 & ~n_8670;
assign n_8672 =  x_1188 & ~n_984;
assign n_8673 = ~n_1021 & ~n_8672;
assign n_8674 =  x_1188 & ~n_8673;
assign n_8675 = ~x_1188 &  n_8673;
assign n_8676 = ~n_8674 & ~n_8675;
assign n_8677 =  x_1187 & ~n_984;
assign n_8678 = ~n_1027 & ~n_8677;
assign n_8679 =  x_1187 & ~n_8678;
assign n_8680 = ~x_1187 &  n_8678;
assign n_8681 = ~n_8679 & ~n_8680;
assign n_8682 =  x_1186 & ~n_984;
assign n_8683 = ~n_1033 & ~n_8682;
assign n_8684 =  x_1186 & ~n_8683;
assign n_8685 = ~x_1186 &  n_8683;
assign n_8686 = ~n_8684 & ~n_8685;
assign n_8687 =  x_1185 & ~n_984;
assign n_8688 = ~n_1039 & ~n_8687;
assign n_8689 =  x_1185 & ~n_8688;
assign n_8690 = ~x_1185 &  n_8688;
assign n_8691 = ~n_8689 & ~n_8690;
assign n_8692 =  x_1184 & ~n_984;
assign n_8693 = ~n_1045 & ~n_8692;
assign n_8694 =  x_1184 & ~n_8693;
assign n_8695 = ~x_1184 &  n_8693;
assign n_8696 = ~n_8694 & ~n_8695;
assign n_8697 =  x_1183 & ~n_984;
assign n_8698 = ~n_1051 & ~n_8697;
assign n_8699 =  x_1183 & ~n_8698;
assign n_8700 = ~x_1183 &  n_8698;
assign n_8701 = ~n_8699 & ~n_8700;
assign n_8702 =  x_1182 & ~n_984;
assign n_8703 = ~n_1057 & ~n_8702;
assign n_8704 =  x_1182 & ~n_8703;
assign n_8705 = ~x_1182 &  n_8703;
assign n_8706 = ~n_8704 & ~n_8705;
assign n_8707 =  x_1181 & ~n_984;
assign n_8708 = ~n_1063 & ~n_8707;
assign n_8709 =  x_1181 & ~n_8708;
assign n_8710 = ~x_1181 &  n_8708;
assign n_8711 = ~n_8709 & ~n_8710;
assign n_8712 =  x_1180 & ~n_984;
assign n_8713 = ~n_1069 & ~n_8712;
assign n_8714 =  x_1180 & ~n_8713;
assign n_8715 = ~x_1180 &  n_8713;
assign n_8716 = ~n_8714 & ~n_8715;
assign n_8717 =  x_1179 & ~n_984;
assign n_8718 = ~n_1075 & ~n_8717;
assign n_8719 =  x_1179 & ~n_8718;
assign n_8720 = ~x_1179 &  n_8718;
assign n_8721 = ~n_8719 & ~n_8720;
assign n_8722 =  x_1178 & ~n_984;
assign n_8723 = ~n_1081 & ~n_8722;
assign n_8724 =  x_1178 & ~n_8723;
assign n_8725 = ~x_1178 &  n_8723;
assign n_8726 = ~n_8724 & ~n_8725;
assign n_8727 =  x_1177 & ~n_984;
assign n_8728 = ~n_1087 & ~n_8727;
assign n_8729 =  x_1177 & ~n_8728;
assign n_8730 = ~x_1177 &  n_8728;
assign n_8731 = ~n_8729 & ~n_8730;
assign n_8732 =  x_1176 & ~n_984;
assign n_8733 = ~n_1093 & ~n_8732;
assign n_8734 =  x_1176 & ~n_8733;
assign n_8735 = ~x_1176 &  n_8733;
assign n_8736 = ~n_8734 & ~n_8735;
assign n_8737 =  x_1175 & ~n_984;
assign n_8738 = ~n_1099 & ~n_8737;
assign n_8739 =  x_1175 & ~n_8738;
assign n_8740 = ~x_1175 &  n_8738;
assign n_8741 = ~n_8739 & ~n_8740;
assign n_8742 =  x_1174 & ~n_984;
assign n_8743 = ~n_1105 & ~n_8742;
assign n_8744 =  x_1174 & ~n_8743;
assign n_8745 = ~x_1174 &  n_8743;
assign n_8746 = ~n_8744 & ~n_8745;
assign n_8747 =  x_1173 & ~n_984;
assign n_8748 = ~n_1111 & ~n_8747;
assign n_8749 =  x_1173 & ~n_8748;
assign n_8750 = ~x_1173 &  n_8748;
assign n_8751 = ~n_8749 & ~n_8750;
assign n_8752 =  x_1172 & ~n_984;
assign n_8753 = ~n_1117 & ~n_8752;
assign n_8754 =  x_1172 & ~n_8753;
assign n_8755 = ~x_1172 &  n_8753;
assign n_8756 = ~n_8754 & ~n_8755;
assign n_8757 =  x_1171 & ~n_984;
assign n_8758 = ~n_1123 & ~n_8757;
assign n_8759 =  x_1171 & ~n_8758;
assign n_8760 = ~x_1171 &  n_8758;
assign n_8761 = ~n_8759 & ~n_8760;
assign n_8762 =  x_1170 & ~n_984;
assign n_8763 = ~n_1129 & ~n_8762;
assign n_8764 =  x_1170 & ~n_8763;
assign n_8765 = ~x_1170 &  n_8763;
assign n_8766 = ~n_8764 & ~n_8765;
assign n_8767 =  x_1169 & ~n_984;
assign n_8768 = ~n_1135 & ~n_8767;
assign n_8769 =  x_1169 & ~n_8768;
assign n_8770 = ~x_1169 &  n_8768;
assign n_8771 = ~n_8769 & ~n_8770;
assign n_8772 =  x_1168 & ~n_984;
assign n_8773 = ~n_1141 & ~n_8772;
assign n_8774 =  x_1168 & ~n_8773;
assign n_8775 = ~x_1168 &  n_8773;
assign n_8776 = ~n_8774 & ~n_8775;
assign n_8777 =  x_1167 & ~n_984;
assign n_8778 = ~n_1147 & ~n_8777;
assign n_8779 =  x_1167 & ~n_8778;
assign n_8780 = ~x_1167 &  n_8778;
assign n_8781 = ~n_8779 & ~n_8780;
assign n_8782 =  x_1166 & ~n_984;
assign n_8783 = ~n_1153 & ~n_8782;
assign n_8784 =  x_1166 & ~n_8783;
assign n_8785 = ~x_1166 &  n_8783;
assign n_8786 = ~n_8784 & ~n_8785;
assign n_8787 =  x_1165 & ~n_984;
assign n_8788 = ~n_1159 & ~n_8787;
assign n_8789 =  x_1165 & ~n_8788;
assign n_8790 = ~x_1165 &  n_8788;
assign n_8791 = ~n_8789 & ~n_8790;
assign n_8792 =  x_1164 & ~n_984;
assign n_8793 = ~n_1165 & ~n_8792;
assign n_8794 =  x_1164 & ~n_8793;
assign n_8795 = ~x_1164 &  n_8793;
assign n_8796 = ~n_8794 & ~n_8795;
assign n_8797 =  x_1163 & ~n_984;
assign n_8798 = ~n_1171 & ~n_8797;
assign n_8799 =  x_1163 & ~n_8798;
assign n_8800 = ~x_1163 &  n_8798;
assign n_8801 = ~n_8799 & ~n_8800;
assign n_8802 =  x_39 &  n_4445;
assign n_8803 =  n_1511 &  n_2886;
assign n_8804 = ~n_2101 & ~n_8803;
assign n_8805 = ~n_8802 &  n_8804;
assign n_8806 =  n_586 & ~n_8805;
assign n_8807 =  x_1162 & ~n_8806;
assign n_8808 =  n_586 &  n_8803;
assign n_8809 =  x_202 &  x_1834;
assign n_8810 = ~x_202 & ~x_1834;
assign n_8811 = ~n_8809 & ~n_8810;
assign n_8812 =  n_8808 &  n_8811;
assign n_8813 =  n_586 &  n_1512;
assign n_8814 =  x_2122 &  x_2794;
assign n_8815 = ~x_2122 & ~x_2794;
assign n_8816 = ~n_8814 & ~n_8815;
assign n_8817 =  n_8813 &  n_8816;
assign n_8818 = ~x_39 &  n_586;
assign n_8819 =  n_8818 &  n_2101;
assign n_8820 =  x_682 &  x_2026;
assign n_8821 = ~x_682 & ~x_2026;
assign n_8822 = ~n_8820 & ~n_8821;
assign n_8823 =  n_8819 &  n_8822;
assign n_8824 =  n_587 &  n_4445;
assign n_8825 =  x_1642 &  n_8824;
assign n_8826 = ~n_8823 & ~n_8825;
assign n_8827 = ~n_8817 &  n_8826;
assign n_8828 = ~n_8812 &  n_8827;
assign n_8829 = ~n_8807 &  n_8828;
assign n_8830 =  x_1162 & ~n_8829;
assign n_8831 = ~x_1162 &  n_8829;
assign n_8832 = ~n_8830 & ~n_8831;
assign n_8833 =  x_1161 & ~n_8806;
assign n_8834 = ~x_1833 & ~x_1834;
assign n_8835 =  x_1833 &  x_1834;
assign n_8836 = ~n_8834 & ~n_8835;
assign n_8837 =  x_201 &  n_8836;
assign n_8838 = ~x_201 & ~n_8836;
assign n_8839 = ~n_8837 & ~n_8838;
assign n_8840 = ~n_8809 & ~n_8839;
assign n_8841 =  n_8809 &  n_8839;
assign n_8842 =  n_8808 & ~n_8841;
assign n_8843 = ~n_8840 &  n_8842;
assign n_8844 = ~x_1641 & ~x_1642;
assign n_8845 =  x_1641 &  x_1642;
assign n_8846 = ~n_8844 & ~n_8845;
assign n_8847 =  n_8824 &  n_8846;
assign n_8848 = ~n_8843 & ~n_8847;
assign n_8849 = ~x_2025 & ~x_2026;
assign n_8850 =  x_2025 &  x_2026;
assign n_8851 = ~n_8849 & ~n_8850;
assign n_8852 =  x_681 &  n_8851;
assign n_8853 = ~x_681 & ~n_8851;
assign n_8854 = ~n_8852 & ~n_8853;
assign n_8855 = ~n_8820 & ~n_8854;
assign n_8856 =  n_8820 &  n_8854;
assign n_8857 =  n_8819 & ~n_8856;
assign n_8858 = ~n_8855 &  n_8857;
assign n_8859 = ~x_2793 & ~x_2794;
assign n_8860 =  x_2793 &  x_2794;
assign n_8861 = ~n_8859 & ~n_8860;
assign n_8862 =  x_2121 &  n_8861;
assign n_8863 = ~x_2121 & ~n_8861;
assign n_8864 = ~n_8862 & ~n_8863;
assign n_8865 =  n_8814 &  n_8864;
assign n_8866 = ~n_8814 & ~n_8864;
assign n_8867 =  n_8813 & ~n_8866;
assign n_8868 = ~n_8865 &  n_8867;
assign n_8869 = ~n_8858 & ~n_8868;
assign n_8870 =  n_8848 &  n_8869;
assign n_8871 = ~n_8833 &  n_8870;
assign n_8872 =  x_1161 & ~n_8871;
assign n_8873 = ~x_1161 &  n_8871;
assign n_8874 = ~n_8872 & ~n_8873;
assign n_8875 = ~x_1832 &  n_8834;
assign n_8876 =  x_1832 & ~n_8834;
assign n_8877 = ~n_8875 & ~n_8876;
assign n_8878 = ~x_201 &  x_1833;
assign n_8879 =  n_8809 & ~n_8878;
assign n_8880 = ~n_8879 & ~n_8837;
assign n_8881 =  n_8877 & ~n_8880;
assign n_8882 = ~n_8877 &  n_8880;
assign n_8883 = ~n_8881 & ~n_8882;
assign n_8884 = ~x_200 & ~n_8883;
assign n_8885 =  x_200 & ~n_8882;
assign n_8886 = ~n_8881 &  n_8885;
assign n_8887 =  n_8808 & ~n_8886;
assign n_8888 = ~n_8884 &  n_8887;
assign n_8889 =  x_1160 & ~n_8806;
assign n_8890 = ~x_1640 &  n_8844;
assign n_8891 =  x_1640 & ~n_8844;
assign n_8892 = ~n_8890 & ~n_8891;
assign n_8893 =  n_8824 &  n_8892;
assign n_8894 = ~n_8889 & ~n_8893;
assign n_8895 = ~n_8888 &  n_8894;
assign n_8896 = ~x_2792 &  n_8859;
assign n_8897 =  x_2792 & ~n_8859;
assign n_8898 = ~n_8896 & ~n_8897;
assign n_8899 = ~x_2121 &  x_2793;
assign n_8900 =  n_8814 & ~n_8899;
assign n_8901 = ~n_8900 & ~n_8862;
assign n_8902 =  n_8898 & ~n_8901;
assign n_8903 = ~n_8898 &  n_8901;
assign n_8904 = ~n_8902 & ~n_8903;
assign n_8905 = ~x_2120 & ~n_8904;
assign n_8906 =  x_2120 & ~n_8903;
assign n_8907 = ~n_8902 &  n_8906;
assign n_8908 =  n_8813 & ~n_8907;
assign n_8909 = ~n_8905 &  n_8908;
assign n_8910 = ~x_2024 &  n_8849;
assign n_8911 =  x_2024 & ~n_8849;
assign n_8912 = ~n_8910 & ~n_8911;
assign n_8913 = ~x_681 &  x_2025;
assign n_8914 =  n_8820 & ~n_8913;
assign n_8915 = ~n_8914 & ~n_8852;
assign n_8916 =  n_8912 & ~n_8915;
assign n_8917 = ~n_8912 &  n_8915;
assign n_8918 = ~n_8916 & ~n_8917;
assign n_8919 =  x_680 &  n_8918;
assign n_8920 = ~x_680 & ~n_8918;
assign n_8921 =  n_8819 & ~n_8920;
assign n_8922 = ~n_8919 &  n_8921;
assign n_8923 = ~n_8909 & ~n_8922;
assign n_8924 =  n_8895 &  n_8923;
assign n_8925 =  x_1160 & ~n_8924;
assign n_8926 = ~x_1160 &  n_8924;
assign n_8927 = ~n_8925 & ~n_8926;
assign n_8928 = ~x_2791 &  n_8896;
assign n_8929 =  x_2791 & ~n_8896;
assign n_8930 = ~n_8928 & ~n_8929;
assign n_8931 = ~n_8902 & ~n_8906;
assign n_8932 =  n_8930 & ~n_8931;
assign n_8933 = ~n_8930 &  n_8931;
assign n_8934 = ~n_8932 & ~n_8933;
assign n_8935 =  x_2119 &  n_8934;
assign n_8936 = ~x_2119 & ~n_8934;
assign n_8937 =  n_8813 & ~n_8936;
assign n_8938 = ~n_8935 &  n_8937;
assign n_8939 =  x_1159 & ~n_8806;
assign n_8940 = ~x_1639 &  n_8890;
assign n_8941 =  x_1639 & ~n_8890;
assign n_8942 = ~n_8940 & ~n_8941;
assign n_8943 =  n_8824 &  n_8942;
assign n_8944 = ~n_8939 & ~n_8943;
assign n_8945 = ~n_8938 &  n_8944;
assign n_8946 = ~x_1831 &  n_8875;
assign n_8947 =  x_1831 & ~n_8875;
assign n_8948 = ~n_8946 & ~n_8947;
assign n_8949 = ~n_8881 & ~n_8885;
assign n_8950 =  n_8948 & ~n_8949;
assign n_8951 = ~n_8948 &  n_8949;
assign n_8952 = ~n_8950 & ~n_8951;
assign n_8953 = ~x_199 & ~n_8952;
assign n_8954 =  x_199 & ~n_8951;
assign n_8955 = ~n_8950 &  n_8954;
assign n_8956 =  n_8808 & ~n_8955;
assign n_8957 = ~n_8953 &  n_8956;
assign n_8958 = ~x_2023 &  n_8910;
assign n_8959 =  x_2023 & ~n_8910;
assign n_8960 = ~n_8958 & ~n_8959;
assign n_8961 =  x_680 & ~n_8917;
assign n_8962 = ~n_8916 & ~n_8961;
assign n_8963 =  n_8960 & ~n_8962;
assign n_8964 = ~n_8960 &  n_8962;
assign n_8965 = ~n_8963 & ~n_8964;
assign n_8966 = ~x_679 & ~n_8965;
assign n_8967 =  x_679 & ~n_8964;
assign n_8968 = ~n_8963 &  n_8967;
assign n_8969 =  n_8819 & ~n_8968;
assign n_8970 = ~n_8966 &  n_8969;
assign n_8971 = ~n_8957 & ~n_8970;
assign n_8972 =  n_8945 &  n_8971;
assign n_8973 =  x_1159 & ~n_8972;
assign n_8974 = ~x_1159 &  n_8972;
assign n_8975 = ~n_8973 & ~n_8974;
assign n_8976 = ~x_2790 &  n_8928;
assign n_8977 =  x_2790 & ~n_8928;
assign n_8978 = ~n_8976 & ~n_8977;
assign n_8979 =  x_2119 & ~n_8933;
assign n_8980 = ~n_8932 & ~n_8979;
assign n_8981 =  n_8978 & ~n_8980;
assign n_8982 = ~n_8978 &  n_8980;
assign n_8983 = ~n_8981 & ~n_8982;
assign n_8984 =  x_2118 &  n_8983;
assign n_8985 = ~x_2118 & ~n_8983;
assign n_8986 =  n_8813 & ~n_8985;
assign n_8987 = ~n_8984 &  n_8986;
assign n_8988 =  x_1158 & ~n_8806;
assign n_8989 =  x_1638 & ~n_8940;
assign n_8990 = ~x_1638 &  n_8940;
assign n_8991 =  n_8824 & ~n_8990;
assign n_8992 = ~n_8989 &  n_8991;
assign n_8993 = ~n_8988 & ~n_8992;
assign n_8994 = ~n_8987 &  n_8993;
assign n_8995 = ~x_1830 &  n_8946;
assign n_8996 =  x_1830 & ~n_8946;
assign n_8997 = ~n_8995 & ~n_8996;
assign n_8998 = ~n_8950 & ~n_8954;
assign n_8999 =  n_8997 & ~n_8998;
assign n_9000 = ~n_8997 &  n_8998;
assign n_9001 = ~n_8999 & ~n_9000;
assign n_9002 = ~x_198 & ~n_9001;
assign n_9003 =  x_198 & ~n_9000;
assign n_9004 = ~n_8999 &  n_9003;
assign n_9005 =  n_8808 & ~n_9004;
assign n_9006 = ~n_9002 &  n_9005;
assign n_9007 = ~x_2022 &  n_8958;
assign n_9008 =  x_2022 & ~n_8958;
assign n_9009 = ~n_9007 & ~n_9008;
assign n_9010 = ~n_8963 & ~n_8967;
assign n_9011 =  n_9009 & ~n_9010;
assign n_9012 = ~n_9009 &  n_9010;
assign n_9013 = ~n_9011 & ~n_9012;
assign n_9014 = ~x_678 & ~n_9013;
assign n_9015 =  x_678 & ~n_9012;
assign n_9016 = ~n_9011 &  n_9015;
assign n_9017 =  n_8819 & ~n_9016;
assign n_9018 = ~n_9014 &  n_9017;
assign n_9019 = ~n_9006 & ~n_9018;
assign n_9020 =  n_8994 &  n_9019;
assign n_9021 =  x_1158 & ~n_9020;
assign n_9022 = ~x_1158 &  n_9020;
assign n_9023 = ~n_9021 & ~n_9022;
assign n_9024 = ~x_2789 &  n_8976;
assign n_9025 =  x_2789 & ~n_8976;
assign n_9026 = ~n_9024 & ~n_9025;
assign n_9027 =  x_2118 & ~n_8982;
assign n_9028 = ~n_8981 & ~n_9027;
assign n_9029 =  n_9026 & ~n_9028;
assign n_9030 = ~n_9026 &  n_9028;
assign n_9031 = ~n_9029 & ~n_9030;
assign n_9032 =  x_2117 &  n_9031;
assign n_9033 = ~x_2117 & ~n_9031;
assign n_9034 =  n_8813 & ~n_9033;
assign n_9035 = ~n_9032 &  n_9034;
assign n_9036 =  x_1157 & ~n_8806;
assign n_9037 =  x_1637 & ~n_8990;
assign n_9038 = ~x_1637 &  n_8990;
assign n_9039 =  n_8824 & ~n_9038;
assign n_9040 = ~n_9037 &  n_9039;
assign n_9041 = ~n_9036 & ~n_9040;
assign n_9042 = ~n_9035 &  n_9041;
assign n_9043 = ~x_1829 &  n_8995;
assign n_9044 =  x_1829 & ~n_8995;
assign n_9045 = ~n_9043 & ~n_9044;
assign n_9046 = ~n_8999 & ~n_9003;
assign n_9047 =  n_9045 & ~n_9046;
assign n_9048 = ~n_9045 &  n_9046;
assign n_9049 = ~n_9047 & ~n_9048;
assign n_9050 = ~x_197 & ~n_9049;
assign n_9051 =  x_197 & ~n_9048;
assign n_9052 = ~n_9047 &  n_9051;
assign n_9053 =  n_8808 & ~n_9052;
assign n_9054 = ~n_9050 &  n_9053;
assign n_9055 = ~x_2021 &  n_9007;
assign n_9056 =  x_2021 & ~n_9007;
assign n_9057 = ~n_9055 & ~n_9056;
assign n_9058 = ~n_9011 & ~n_9015;
assign n_9059 =  n_9057 & ~n_9058;
assign n_9060 = ~n_9057 &  n_9058;
assign n_9061 = ~n_9059 & ~n_9060;
assign n_9062 = ~x_677 & ~n_9061;
assign n_9063 =  x_677 & ~n_9060;
assign n_9064 = ~n_9059 &  n_9063;
assign n_9065 =  n_8819 & ~n_9064;
assign n_9066 = ~n_9062 &  n_9065;
assign n_9067 = ~n_9054 & ~n_9066;
assign n_9068 =  n_9042 &  n_9067;
assign n_9069 =  x_1157 & ~n_9068;
assign n_9070 = ~x_1157 &  n_9068;
assign n_9071 = ~n_9069 & ~n_9070;
assign n_9072 = ~x_2788 &  n_9024;
assign n_9073 =  x_2788 & ~n_9024;
assign n_9074 = ~n_9072 & ~n_9073;
assign n_9075 =  x_2117 & ~n_9030;
assign n_9076 = ~n_9029 & ~n_9075;
assign n_9077 =  n_9074 & ~n_9076;
assign n_9078 = ~n_9074 &  n_9076;
assign n_9079 = ~n_9077 & ~n_9078;
assign n_9080 =  x_2116 &  n_9079;
assign n_9081 = ~x_2116 & ~n_9079;
assign n_9082 =  n_8813 & ~n_9081;
assign n_9083 = ~n_9080 &  n_9082;
assign n_9084 =  x_1156 & ~n_8806;
assign n_9085 =  x_1636 & ~n_9038;
assign n_9086 = ~x_1636 &  n_9038;
assign n_9087 =  n_8824 & ~n_9086;
assign n_9088 = ~n_9085 &  n_9087;
assign n_9089 = ~n_9084 & ~n_9088;
assign n_9090 = ~n_9083 &  n_9089;
assign n_9091 = ~x_1828 &  n_9043;
assign n_9092 =  x_1828 & ~n_9043;
assign n_9093 = ~n_9091 & ~n_9092;
assign n_9094 = ~n_9047 & ~n_9051;
assign n_9095 =  n_9093 & ~n_9094;
assign n_9096 = ~n_9093 &  n_9094;
assign n_9097 = ~n_9095 & ~n_9096;
assign n_9098 = ~x_196 & ~n_9097;
assign n_9099 =  x_196 & ~n_9096;
assign n_9100 = ~n_9095 &  n_9099;
assign n_9101 =  n_8808 & ~n_9100;
assign n_9102 = ~n_9098 &  n_9101;
assign n_9103 = ~x_2020 &  n_9055;
assign n_9104 =  x_2020 & ~n_9055;
assign n_9105 = ~n_9103 & ~n_9104;
assign n_9106 = ~n_9059 & ~n_9063;
assign n_9107 =  n_9105 & ~n_9106;
assign n_9108 = ~n_9105 &  n_9106;
assign n_9109 = ~n_9107 & ~n_9108;
assign n_9110 = ~x_676 & ~n_9109;
assign n_9111 =  x_676 & ~n_9108;
assign n_9112 = ~n_9107 &  n_9111;
assign n_9113 =  n_8819 & ~n_9112;
assign n_9114 = ~n_9110 &  n_9113;
assign n_9115 = ~n_9102 & ~n_9114;
assign n_9116 =  n_9090 &  n_9115;
assign n_9117 =  x_1156 & ~n_9116;
assign n_9118 = ~x_1156 &  n_9116;
assign n_9119 = ~n_9117 & ~n_9118;
assign n_9120 = ~x_2787 &  n_9072;
assign n_9121 =  x_2787 & ~n_9072;
assign n_9122 = ~n_9120 & ~n_9121;
assign n_9123 =  x_2116 & ~n_9078;
assign n_9124 = ~n_9077 & ~n_9123;
assign n_9125 =  n_9122 & ~n_9124;
assign n_9126 = ~n_9122 &  n_9124;
assign n_9127 = ~n_9125 & ~n_9126;
assign n_9128 =  x_2115 &  n_9127;
assign n_9129 = ~x_2115 & ~n_9127;
assign n_9130 =  n_8813 & ~n_9129;
assign n_9131 = ~n_9128 &  n_9130;
assign n_9132 =  x_1155 & ~n_8806;
assign n_9133 =  x_1635 & ~n_9086;
assign n_9134 = ~x_1635 &  n_9086;
assign n_9135 =  n_8824 & ~n_9134;
assign n_9136 = ~n_9133 &  n_9135;
assign n_9137 = ~n_9132 & ~n_9136;
assign n_9138 = ~n_9131 &  n_9137;
assign n_9139 = ~x_1827 &  n_9091;
assign n_9140 =  x_1827 & ~n_9091;
assign n_9141 = ~n_9139 & ~n_9140;
assign n_9142 = ~n_9095 & ~n_9099;
assign n_9143 =  n_9141 & ~n_9142;
assign n_9144 = ~n_9141 &  n_9142;
assign n_9145 = ~n_9143 & ~n_9144;
assign n_9146 = ~x_195 & ~n_9145;
assign n_9147 =  x_195 & ~n_9144;
assign n_9148 = ~n_9143 &  n_9147;
assign n_9149 =  n_8808 & ~n_9148;
assign n_9150 = ~n_9146 &  n_9149;
assign n_9151 = ~x_2019 &  n_9103;
assign n_9152 =  x_2019 & ~n_9103;
assign n_9153 = ~n_9151 & ~n_9152;
assign n_9154 = ~n_9107 & ~n_9111;
assign n_9155 =  n_9153 & ~n_9154;
assign n_9156 = ~n_9153 &  n_9154;
assign n_9157 = ~n_9155 & ~n_9156;
assign n_9158 = ~x_675 & ~n_9157;
assign n_9159 =  x_675 & ~n_9156;
assign n_9160 = ~n_9155 &  n_9159;
assign n_9161 =  n_8819 & ~n_9160;
assign n_9162 = ~n_9158 &  n_9161;
assign n_9163 = ~n_9150 & ~n_9162;
assign n_9164 =  n_9138 &  n_9163;
assign n_9165 =  x_1155 & ~n_9164;
assign n_9166 = ~x_1155 &  n_9164;
assign n_9167 = ~n_9165 & ~n_9166;
assign n_9168 = ~x_2786 &  n_9120;
assign n_9169 =  x_2786 & ~n_9120;
assign n_9170 = ~n_9168 & ~n_9169;
assign n_9171 =  x_2115 & ~n_9126;
assign n_9172 = ~n_9125 & ~n_9171;
assign n_9173 =  n_9170 & ~n_9172;
assign n_9174 = ~n_9170 &  n_9172;
assign n_9175 = ~n_9173 & ~n_9174;
assign n_9176 =  x_2114 &  n_9175;
assign n_9177 = ~x_2114 & ~n_9175;
assign n_9178 =  n_8813 & ~n_9177;
assign n_9179 = ~n_9176 &  n_9178;
assign n_9180 =  x_1154 & ~n_8806;
assign n_9181 =  x_1634 & ~n_9134;
assign n_9182 = ~x_1634 &  n_9134;
assign n_9183 =  n_8824 & ~n_9182;
assign n_9184 = ~n_9181 &  n_9183;
assign n_9185 = ~n_9180 & ~n_9184;
assign n_9186 = ~n_9179 &  n_9185;
assign n_9187 = ~x_1826 &  n_9139;
assign n_9188 =  x_1826 & ~n_9139;
assign n_9189 = ~n_9187 & ~n_9188;
assign n_9190 = ~n_9143 & ~n_9147;
assign n_9191 =  n_9189 & ~n_9190;
assign n_9192 = ~n_9189 &  n_9190;
assign n_9193 = ~n_9191 & ~n_9192;
assign n_9194 = ~x_194 & ~n_9193;
assign n_9195 =  x_194 & ~n_9192;
assign n_9196 = ~n_9191 &  n_9195;
assign n_9197 =  n_8808 & ~n_9196;
assign n_9198 = ~n_9194 &  n_9197;
assign n_9199 = ~x_2018 &  n_9151;
assign n_9200 =  x_2018 & ~n_9151;
assign n_9201 = ~n_9199 & ~n_9200;
assign n_9202 = ~n_9155 & ~n_9159;
assign n_9203 =  n_9201 & ~n_9202;
assign n_9204 = ~n_9201 &  n_9202;
assign n_9205 = ~n_9203 & ~n_9204;
assign n_9206 = ~x_674 & ~n_9205;
assign n_9207 =  x_674 & ~n_9204;
assign n_9208 = ~n_9203 &  n_9207;
assign n_9209 =  n_8819 & ~n_9208;
assign n_9210 = ~n_9206 &  n_9209;
assign n_9211 = ~n_9198 & ~n_9210;
assign n_9212 =  n_9186 &  n_9211;
assign n_9213 =  x_1154 & ~n_9212;
assign n_9214 = ~x_1154 &  n_9212;
assign n_9215 = ~n_9213 & ~n_9214;
assign n_9216 = ~x_2785 &  n_9168;
assign n_9217 =  x_2785 & ~n_9168;
assign n_9218 = ~n_9216 & ~n_9217;
assign n_9219 =  x_2114 & ~n_9174;
assign n_9220 = ~n_9173 & ~n_9219;
assign n_9221 =  n_9218 & ~n_9220;
assign n_9222 = ~n_9218 &  n_9220;
assign n_9223 = ~n_9221 & ~n_9222;
assign n_9224 =  x_2113 &  n_9223;
assign n_9225 = ~x_2113 & ~n_9223;
assign n_9226 =  n_8813 & ~n_9225;
assign n_9227 = ~n_9224 &  n_9226;
assign n_9228 =  x_1153 & ~n_8806;
assign n_9229 =  x_1633 & ~n_9182;
assign n_9230 = ~x_1633 &  n_9182;
assign n_9231 =  n_8824 & ~n_9230;
assign n_9232 = ~n_9229 &  n_9231;
assign n_9233 = ~n_9228 & ~n_9232;
assign n_9234 = ~n_9227 &  n_9233;
assign n_9235 = ~x_1825 &  n_9187;
assign n_9236 =  x_1825 & ~n_9187;
assign n_9237 = ~n_9235 & ~n_9236;
assign n_9238 = ~n_9191 & ~n_9195;
assign n_9239 =  n_9237 & ~n_9238;
assign n_9240 = ~n_9237 &  n_9238;
assign n_9241 = ~n_9239 & ~n_9240;
assign n_9242 = ~x_193 & ~n_9241;
assign n_9243 =  x_193 & ~n_9240;
assign n_9244 = ~n_9239 &  n_9243;
assign n_9245 =  n_8808 & ~n_9244;
assign n_9246 = ~n_9242 &  n_9245;
assign n_9247 = ~x_2017 &  n_9199;
assign n_9248 =  x_2017 & ~n_9199;
assign n_9249 = ~n_9247 & ~n_9248;
assign n_9250 = ~n_9203 & ~n_9207;
assign n_9251 =  n_9249 & ~n_9250;
assign n_9252 = ~n_9249 &  n_9250;
assign n_9253 = ~n_9251 & ~n_9252;
assign n_9254 = ~x_673 & ~n_9253;
assign n_9255 =  x_673 & ~n_9252;
assign n_9256 = ~n_9251 &  n_9255;
assign n_9257 =  n_8819 & ~n_9256;
assign n_9258 = ~n_9254 &  n_9257;
assign n_9259 = ~n_9246 & ~n_9258;
assign n_9260 =  n_9234 &  n_9259;
assign n_9261 =  x_1153 & ~n_9260;
assign n_9262 = ~x_1153 &  n_9260;
assign n_9263 = ~n_9261 & ~n_9262;
assign n_9264 = ~x_2784 &  n_9216;
assign n_9265 =  x_2784 & ~n_9216;
assign n_9266 = ~n_9264 & ~n_9265;
assign n_9267 =  x_2113 & ~n_9222;
assign n_9268 = ~n_9221 & ~n_9267;
assign n_9269 =  n_9266 & ~n_9268;
assign n_9270 = ~n_9266 &  n_9268;
assign n_9271 = ~n_9269 & ~n_9270;
assign n_9272 =  x_2112 &  n_9271;
assign n_9273 = ~x_2112 & ~n_9271;
assign n_9274 =  n_8813 & ~n_9273;
assign n_9275 = ~n_9272 &  n_9274;
assign n_9276 =  x_1152 & ~n_8806;
assign n_9277 =  x_1632 & ~n_9230;
assign n_9278 = ~x_1632 &  n_9230;
assign n_9279 =  n_8824 & ~n_9278;
assign n_9280 = ~n_9277 &  n_9279;
assign n_9281 = ~n_9276 & ~n_9280;
assign n_9282 = ~n_9275 &  n_9281;
assign n_9283 = ~x_1824 &  n_9235;
assign n_9284 =  x_1824 & ~n_9235;
assign n_9285 = ~n_9283 & ~n_9284;
assign n_9286 = ~n_9239 & ~n_9243;
assign n_9287 =  n_9285 & ~n_9286;
assign n_9288 = ~n_9285 &  n_9286;
assign n_9289 = ~n_9287 & ~n_9288;
assign n_9290 = ~x_192 & ~n_9289;
assign n_9291 =  x_192 & ~n_9288;
assign n_9292 = ~n_9287 &  n_9291;
assign n_9293 =  n_8808 & ~n_9292;
assign n_9294 = ~n_9290 &  n_9293;
assign n_9295 = ~x_2016 &  n_9247;
assign n_9296 =  x_2016 & ~n_9247;
assign n_9297 = ~n_9295 & ~n_9296;
assign n_9298 = ~n_9251 & ~n_9255;
assign n_9299 =  n_9297 & ~n_9298;
assign n_9300 = ~n_9297 &  n_9298;
assign n_9301 = ~n_9299 & ~n_9300;
assign n_9302 = ~x_672 & ~n_9301;
assign n_9303 =  x_672 & ~n_9300;
assign n_9304 = ~n_9299 &  n_9303;
assign n_9305 =  n_8819 & ~n_9304;
assign n_9306 = ~n_9302 &  n_9305;
assign n_9307 = ~n_9294 & ~n_9306;
assign n_9308 =  n_9282 &  n_9307;
assign n_9309 =  x_1152 & ~n_9308;
assign n_9310 = ~x_1152 &  n_9308;
assign n_9311 = ~n_9309 & ~n_9310;
assign n_9312 = ~x_2783 &  n_9264;
assign n_9313 =  x_2783 & ~n_9264;
assign n_9314 = ~n_9312 & ~n_9313;
assign n_9315 =  x_2112 & ~n_9270;
assign n_9316 = ~n_9269 & ~n_9315;
assign n_9317 =  n_9314 & ~n_9316;
assign n_9318 = ~n_9314 &  n_9316;
assign n_9319 = ~n_9317 & ~n_9318;
assign n_9320 =  x_2111 &  n_9319;
assign n_9321 = ~x_2111 & ~n_9319;
assign n_9322 =  n_8813 & ~n_9321;
assign n_9323 = ~n_9320 &  n_9322;
assign n_9324 =  x_1151 & ~n_8806;
assign n_9325 =  x_1631 & ~n_9278;
assign n_9326 = ~x_1631 &  n_9278;
assign n_9327 =  n_8824 & ~n_9326;
assign n_9328 = ~n_9325 &  n_9327;
assign n_9329 = ~n_9324 & ~n_9328;
assign n_9330 = ~n_9323 &  n_9329;
assign n_9331 = ~x_1823 &  n_9283;
assign n_9332 =  x_1823 & ~n_9283;
assign n_9333 = ~n_9331 & ~n_9332;
assign n_9334 = ~n_9287 & ~n_9291;
assign n_9335 =  n_9333 & ~n_9334;
assign n_9336 = ~n_9333 &  n_9334;
assign n_9337 = ~n_9335 & ~n_9336;
assign n_9338 = ~x_191 & ~n_9337;
assign n_9339 =  x_191 & ~n_9336;
assign n_9340 = ~n_9335 &  n_9339;
assign n_9341 =  n_8808 & ~n_9340;
assign n_9342 = ~n_9338 &  n_9341;
assign n_9343 = ~x_2015 &  n_9295;
assign n_9344 =  x_2015 & ~n_9295;
assign n_9345 = ~n_9343 & ~n_9344;
assign n_9346 = ~n_9299 & ~n_9303;
assign n_9347 =  n_9345 & ~n_9346;
assign n_9348 = ~n_9345 &  n_9346;
assign n_9349 = ~n_9347 & ~n_9348;
assign n_9350 = ~x_671 & ~n_9349;
assign n_9351 =  x_671 & ~n_9348;
assign n_9352 = ~n_9347 &  n_9351;
assign n_9353 =  n_8819 & ~n_9352;
assign n_9354 = ~n_9350 &  n_9353;
assign n_9355 = ~n_9342 & ~n_9354;
assign n_9356 =  n_9330 &  n_9355;
assign n_9357 =  x_1151 & ~n_9356;
assign n_9358 = ~x_1151 &  n_9356;
assign n_9359 = ~n_9357 & ~n_9358;
assign n_9360 = ~x_2782 &  n_9312;
assign n_9361 =  x_2782 & ~n_9312;
assign n_9362 = ~n_9360 & ~n_9361;
assign n_9363 =  x_2111 & ~n_9318;
assign n_9364 = ~n_9317 & ~n_9363;
assign n_9365 =  n_9362 & ~n_9364;
assign n_9366 = ~n_9362 &  n_9364;
assign n_9367 = ~n_9365 & ~n_9366;
assign n_9368 =  x_2110 &  n_9367;
assign n_9369 = ~x_2110 & ~n_9367;
assign n_9370 =  n_8813 & ~n_9369;
assign n_9371 = ~n_9368 &  n_9370;
assign n_9372 =  x_1150 & ~n_8806;
assign n_9373 =  x_1630 & ~n_9326;
assign n_9374 = ~x_1630 &  n_9326;
assign n_9375 =  n_8824 & ~n_9374;
assign n_9376 = ~n_9373 &  n_9375;
assign n_9377 = ~n_9372 & ~n_9376;
assign n_9378 = ~n_9371 &  n_9377;
assign n_9379 = ~x_1822 &  n_9331;
assign n_9380 =  x_1822 & ~n_9331;
assign n_9381 = ~n_9379 & ~n_9380;
assign n_9382 = ~n_9335 & ~n_9339;
assign n_9383 =  n_9381 & ~n_9382;
assign n_9384 = ~n_9381 &  n_9382;
assign n_9385 = ~n_9383 & ~n_9384;
assign n_9386 = ~x_190 & ~n_9385;
assign n_9387 =  x_190 & ~n_9384;
assign n_9388 = ~n_9383 &  n_9387;
assign n_9389 =  n_8808 & ~n_9388;
assign n_9390 = ~n_9386 &  n_9389;
assign n_9391 = ~x_2014 &  n_9343;
assign n_9392 =  x_2014 & ~n_9343;
assign n_9393 = ~n_9391 & ~n_9392;
assign n_9394 = ~n_9347 & ~n_9351;
assign n_9395 =  n_9393 & ~n_9394;
assign n_9396 = ~n_9393 &  n_9394;
assign n_9397 = ~n_9395 & ~n_9396;
assign n_9398 = ~x_670 & ~n_9397;
assign n_9399 =  x_670 & ~n_9396;
assign n_9400 = ~n_9395 &  n_9399;
assign n_9401 =  n_8819 & ~n_9400;
assign n_9402 = ~n_9398 &  n_9401;
assign n_9403 = ~n_9390 & ~n_9402;
assign n_9404 =  n_9378 &  n_9403;
assign n_9405 =  x_1150 & ~n_9404;
assign n_9406 = ~x_1150 &  n_9404;
assign n_9407 = ~n_9405 & ~n_9406;
assign n_9408 = ~x_2781 &  n_9360;
assign n_9409 =  x_2781 & ~n_9360;
assign n_9410 = ~n_9408 & ~n_9409;
assign n_9411 =  x_2110 & ~n_9366;
assign n_9412 = ~n_9365 & ~n_9411;
assign n_9413 =  n_9410 & ~n_9412;
assign n_9414 = ~n_9410 &  n_9412;
assign n_9415 = ~n_9413 & ~n_9414;
assign n_9416 =  x_2109 &  n_9415;
assign n_9417 = ~x_2109 & ~n_9415;
assign n_9418 =  n_8813 & ~n_9417;
assign n_9419 = ~n_9416 &  n_9418;
assign n_9420 =  x_1149 & ~n_8806;
assign n_9421 =  x_1629 & ~n_9374;
assign n_9422 = ~x_1629 &  n_9374;
assign n_9423 =  n_8824 & ~n_9422;
assign n_9424 = ~n_9421 &  n_9423;
assign n_9425 = ~n_9420 & ~n_9424;
assign n_9426 = ~n_9419 &  n_9425;
assign n_9427 = ~x_1821 &  n_9379;
assign n_9428 =  x_1821 & ~n_9379;
assign n_9429 = ~n_9427 & ~n_9428;
assign n_9430 = ~n_9383 & ~n_9387;
assign n_9431 =  n_9429 & ~n_9430;
assign n_9432 = ~n_9429 &  n_9430;
assign n_9433 = ~n_9431 & ~n_9432;
assign n_9434 = ~x_189 & ~n_9433;
assign n_9435 =  x_189 & ~n_9432;
assign n_9436 = ~n_9431 &  n_9435;
assign n_9437 =  n_8808 & ~n_9436;
assign n_9438 = ~n_9434 &  n_9437;
assign n_9439 = ~x_2013 &  n_9391;
assign n_9440 =  x_2013 & ~n_9391;
assign n_9441 = ~n_9439 & ~n_9440;
assign n_9442 = ~n_9395 & ~n_9399;
assign n_9443 =  n_9441 & ~n_9442;
assign n_9444 = ~n_9441 &  n_9442;
assign n_9445 = ~n_9443 & ~n_9444;
assign n_9446 = ~x_669 & ~n_9445;
assign n_9447 =  x_669 & ~n_9444;
assign n_9448 = ~n_9443 &  n_9447;
assign n_9449 =  n_8819 & ~n_9448;
assign n_9450 = ~n_9446 &  n_9449;
assign n_9451 = ~n_9438 & ~n_9450;
assign n_9452 =  n_9426 &  n_9451;
assign n_9453 =  x_1149 & ~n_9452;
assign n_9454 = ~x_1149 &  n_9452;
assign n_9455 = ~n_9453 & ~n_9454;
assign n_9456 = ~x_2780 &  n_9408;
assign n_9457 =  x_2780 & ~n_9408;
assign n_9458 = ~n_9456 & ~n_9457;
assign n_9459 =  x_2109 & ~n_9414;
assign n_9460 = ~n_9413 & ~n_9459;
assign n_9461 =  n_9458 & ~n_9460;
assign n_9462 = ~n_9458 &  n_9460;
assign n_9463 = ~n_9461 & ~n_9462;
assign n_9464 =  x_2108 &  n_9463;
assign n_9465 = ~x_2108 & ~n_9463;
assign n_9466 =  n_8813 & ~n_9465;
assign n_9467 = ~n_9464 &  n_9466;
assign n_9468 =  x_1148 & ~n_8806;
assign n_9469 =  x_1628 & ~n_9422;
assign n_9470 = ~x_1628 &  n_9422;
assign n_9471 =  n_8824 & ~n_9470;
assign n_9472 = ~n_9469 &  n_9471;
assign n_9473 = ~n_9468 & ~n_9472;
assign n_9474 = ~n_9467 &  n_9473;
assign n_9475 = ~x_1820 &  n_9427;
assign n_9476 =  x_1820 & ~n_9427;
assign n_9477 = ~n_9475 & ~n_9476;
assign n_9478 = ~n_9431 & ~n_9435;
assign n_9479 =  n_9477 & ~n_9478;
assign n_9480 = ~n_9477 &  n_9478;
assign n_9481 = ~n_9479 & ~n_9480;
assign n_9482 = ~x_188 & ~n_9481;
assign n_9483 =  x_188 & ~n_9480;
assign n_9484 = ~n_9479 &  n_9483;
assign n_9485 =  n_8808 & ~n_9484;
assign n_9486 = ~n_9482 &  n_9485;
assign n_9487 = ~x_2012 &  n_9439;
assign n_9488 =  x_2012 & ~n_9439;
assign n_9489 = ~n_9487 & ~n_9488;
assign n_9490 = ~n_9443 & ~n_9447;
assign n_9491 =  n_9489 & ~n_9490;
assign n_9492 = ~n_9489 &  n_9490;
assign n_9493 = ~n_9491 & ~n_9492;
assign n_9494 = ~x_668 & ~n_9493;
assign n_9495 =  x_668 & ~n_9492;
assign n_9496 = ~n_9491 &  n_9495;
assign n_9497 =  n_8819 & ~n_9496;
assign n_9498 = ~n_9494 &  n_9497;
assign n_9499 = ~n_9486 & ~n_9498;
assign n_9500 =  n_9474 &  n_9499;
assign n_9501 =  x_1148 & ~n_9500;
assign n_9502 = ~x_1148 &  n_9500;
assign n_9503 = ~n_9501 & ~n_9502;
assign n_9504 = ~x_2779 &  n_9456;
assign n_9505 =  x_2779 & ~n_9456;
assign n_9506 = ~n_9504 & ~n_9505;
assign n_9507 =  x_2108 & ~n_9462;
assign n_9508 = ~n_9461 & ~n_9507;
assign n_9509 =  n_9506 & ~n_9508;
assign n_9510 = ~n_9506 &  n_9508;
assign n_9511 = ~n_9509 & ~n_9510;
assign n_9512 =  x_2107 &  n_9511;
assign n_9513 = ~x_2107 & ~n_9511;
assign n_9514 =  n_8813 & ~n_9513;
assign n_9515 = ~n_9512 &  n_9514;
assign n_9516 =  x_1147 & ~n_8806;
assign n_9517 =  x_1627 & ~n_9470;
assign n_9518 = ~x_1627 &  n_9470;
assign n_9519 =  n_8824 & ~n_9518;
assign n_9520 = ~n_9517 &  n_9519;
assign n_9521 = ~n_9516 & ~n_9520;
assign n_9522 = ~n_9515 &  n_9521;
assign n_9523 = ~x_1819 &  n_9475;
assign n_9524 =  x_1819 & ~n_9475;
assign n_9525 = ~n_9523 & ~n_9524;
assign n_9526 = ~n_9479 & ~n_9483;
assign n_9527 =  n_9525 & ~n_9526;
assign n_9528 = ~n_9525 &  n_9526;
assign n_9529 = ~n_9527 & ~n_9528;
assign n_9530 = ~x_187 & ~n_9529;
assign n_9531 =  x_187 & ~n_9528;
assign n_9532 = ~n_9527 &  n_9531;
assign n_9533 =  n_8808 & ~n_9532;
assign n_9534 = ~n_9530 &  n_9533;
assign n_9535 = ~x_2011 &  n_9487;
assign n_9536 =  x_2011 & ~n_9487;
assign n_9537 = ~n_9535 & ~n_9536;
assign n_9538 = ~n_9491 & ~n_9495;
assign n_9539 =  n_9537 & ~n_9538;
assign n_9540 = ~n_9537 &  n_9538;
assign n_9541 = ~n_9539 & ~n_9540;
assign n_9542 = ~x_667 & ~n_9541;
assign n_9543 =  x_667 & ~n_9540;
assign n_9544 = ~n_9539 &  n_9543;
assign n_9545 =  n_8819 & ~n_9544;
assign n_9546 = ~n_9542 &  n_9545;
assign n_9547 = ~n_9534 & ~n_9546;
assign n_9548 =  n_9522 &  n_9547;
assign n_9549 =  x_1147 & ~n_9548;
assign n_9550 = ~x_1147 &  n_9548;
assign n_9551 = ~n_9549 & ~n_9550;
assign n_9552 = ~x_2778 &  n_9504;
assign n_9553 =  x_2778 & ~n_9504;
assign n_9554 = ~n_9552 & ~n_9553;
assign n_9555 =  x_2107 & ~n_9510;
assign n_9556 = ~n_9509 & ~n_9555;
assign n_9557 =  n_9554 & ~n_9556;
assign n_9558 = ~n_9554 &  n_9556;
assign n_9559 = ~n_9557 & ~n_9558;
assign n_9560 =  x_2106 &  n_9559;
assign n_9561 = ~x_2106 & ~n_9559;
assign n_9562 =  n_8813 & ~n_9561;
assign n_9563 = ~n_9560 &  n_9562;
assign n_9564 =  x_1146 & ~n_8806;
assign n_9565 =  x_1626 & ~n_9518;
assign n_9566 = ~x_1626 &  n_9518;
assign n_9567 =  n_8824 & ~n_9566;
assign n_9568 = ~n_9565 &  n_9567;
assign n_9569 = ~n_9564 & ~n_9568;
assign n_9570 = ~n_9563 &  n_9569;
assign n_9571 = ~x_1818 &  n_9523;
assign n_9572 =  x_1818 & ~n_9523;
assign n_9573 = ~n_9571 & ~n_9572;
assign n_9574 = ~n_9527 & ~n_9531;
assign n_9575 =  n_9573 & ~n_9574;
assign n_9576 = ~n_9573 &  n_9574;
assign n_9577 = ~n_9575 & ~n_9576;
assign n_9578 = ~x_186 & ~n_9577;
assign n_9579 =  x_186 & ~n_9576;
assign n_9580 = ~n_9575 &  n_9579;
assign n_9581 =  n_8808 & ~n_9580;
assign n_9582 = ~n_9578 &  n_9581;
assign n_9583 = ~x_2010 &  n_9535;
assign n_9584 =  x_2010 & ~n_9535;
assign n_9585 = ~n_9583 & ~n_9584;
assign n_9586 = ~n_9539 & ~n_9543;
assign n_9587 =  n_9585 & ~n_9586;
assign n_9588 = ~n_9585 &  n_9586;
assign n_9589 = ~n_9587 & ~n_9588;
assign n_9590 = ~x_666 & ~n_9589;
assign n_9591 =  x_666 & ~n_9588;
assign n_9592 = ~n_9587 &  n_9591;
assign n_9593 =  n_8819 & ~n_9592;
assign n_9594 = ~n_9590 &  n_9593;
assign n_9595 = ~n_9582 & ~n_9594;
assign n_9596 =  n_9570 &  n_9595;
assign n_9597 =  x_1146 & ~n_9596;
assign n_9598 = ~x_1146 &  n_9596;
assign n_9599 = ~n_9597 & ~n_9598;
assign n_9600 = ~x_2777 &  n_9552;
assign n_9601 =  x_2777 & ~n_9552;
assign n_9602 = ~n_9600 & ~n_9601;
assign n_9603 =  x_2106 & ~n_9558;
assign n_9604 = ~n_9557 & ~n_9603;
assign n_9605 =  n_9602 & ~n_9604;
assign n_9606 = ~n_9602 &  n_9604;
assign n_9607 = ~n_9605 & ~n_9606;
assign n_9608 =  x_2105 &  n_9607;
assign n_9609 = ~x_2105 & ~n_9607;
assign n_9610 =  n_8813 & ~n_9609;
assign n_9611 = ~n_9608 &  n_9610;
assign n_9612 =  x_1145 & ~n_8806;
assign n_9613 =  x_1625 & ~n_9566;
assign n_9614 = ~x_1625 &  n_9566;
assign n_9615 =  n_8824 & ~n_9614;
assign n_9616 = ~n_9613 &  n_9615;
assign n_9617 = ~n_9612 & ~n_9616;
assign n_9618 = ~n_9611 &  n_9617;
assign n_9619 = ~x_1817 &  n_9571;
assign n_9620 =  x_1817 & ~n_9571;
assign n_9621 = ~n_9619 & ~n_9620;
assign n_9622 = ~n_9575 & ~n_9579;
assign n_9623 =  n_9621 & ~n_9622;
assign n_9624 = ~n_9621 &  n_9622;
assign n_9625 = ~n_9623 & ~n_9624;
assign n_9626 = ~x_185 & ~n_9625;
assign n_9627 =  x_185 & ~n_9624;
assign n_9628 = ~n_9623 &  n_9627;
assign n_9629 =  n_8808 & ~n_9628;
assign n_9630 = ~n_9626 &  n_9629;
assign n_9631 = ~x_2009 &  n_9583;
assign n_9632 =  x_2009 & ~n_9583;
assign n_9633 = ~n_9631 & ~n_9632;
assign n_9634 = ~n_9587 & ~n_9591;
assign n_9635 =  n_9633 & ~n_9634;
assign n_9636 = ~n_9633 &  n_9634;
assign n_9637 = ~n_9635 & ~n_9636;
assign n_9638 = ~x_665 & ~n_9637;
assign n_9639 =  x_665 & ~n_9636;
assign n_9640 = ~n_9635 &  n_9639;
assign n_9641 =  n_8819 & ~n_9640;
assign n_9642 = ~n_9638 &  n_9641;
assign n_9643 = ~n_9630 & ~n_9642;
assign n_9644 =  n_9618 &  n_9643;
assign n_9645 =  x_1145 & ~n_9644;
assign n_9646 = ~x_1145 &  n_9644;
assign n_9647 = ~n_9645 & ~n_9646;
assign n_9648 = ~x_2776 &  n_9600;
assign n_9649 =  x_2776 & ~n_9600;
assign n_9650 = ~n_9648 & ~n_9649;
assign n_9651 =  x_2105 & ~n_9606;
assign n_9652 = ~n_9605 & ~n_9651;
assign n_9653 =  n_9650 & ~n_9652;
assign n_9654 = ~n_9650 &  n_9652;
assign n_9655 = ~n_9653 & ~n_9654;
assign n_9656 =  x_2104 &  n_9655;
assign n_9657 = ~x_2104 & ~n_9655;
assign n_9658 =  n_8813 & ~n_9657;
assign n_9659 = ~n_9656 &  n_9658;
assign n_9660 =  x_1144 & ~n_8806;
assign n_9661 =  x_1624 & ~n_9614;
assign n_9662 = ~x_1624 &  n_9614;
assign n_9663 =  n_8824 & ~n_9662;
assign n_9664 = ~n_9661 &  n_9663;
assign n_9665 = ~n_9660 & ~n_9664;
assign n_9666 = ~n_9659 &  n_9665;
assign n_9667 = ~x_1816 &  n_9619;
assign n_9668 =  x_1816 & ~n_9619;
assign n_9669 = ~n_9667 & ~n_9668;
assign n_9670 = ~n_9623 & ~n_9627;
assign n_9671 =  n_9669 & ~n_9670;
assign n_9672 = ~n_9669 &  n_9670;
assign n_9673 = ~n_9671 & ~n_9672;
assign n_9674 = ~x_184 & ~n_9673;
assign n_9675 =  x_184 & ~n_9672;
assign n_9676 = ~n_9671 &  n_9675;
assign n_9677 =  n_8808 & ~n_9676;
assign n_9678 = ~n_9674 &  n_9677;
assign n_9679 = ~x_2008 &  n_9631;
assign n_9680 =  x_2008 & ~n_9631;
assign n_9681 = ~n_9679 & ~n_9680;
assign n_9682 = ~n_9635 & ~n_9639;
assign n_9683 =  n_9681 & ~n_9682;
assign n_9684 = ~n_9681 &  n_9682;
assign n_9685 = ~n_9683 & ~n_9684;
assign n_9686 = ~x_664 & ~n_9685;
assign n_9687 =  x_664 & ~n_9684;
assign n_9688 = ~n_9683 &  n_9687;
assign n_9689 =  n_8819 & ~n_9688;
assign n_9690 = ~n_9686 &  n_9689;
assign n_9691 = ~n_9678 & ~n_9690;
assign n_9692 =  n_9666 &  n_9691;
assign n_9693 =  x_1144 & ~n_9692;
assign n_9694 = ~x_1144 &  n_9692;
assign n_9695 = ~n_9693 & ~n_9694;
assign n_9696 = ~x_2775 &  n_9648;
assign n_9697 =  x_2775 & ~n_9648;
assign n_9698 = ~n_9696 & ~n_9697;
assign n_9699 =  x_2104 & ~n_9654;
assign n_9700 = ~n_9653 & ~n_9699;
assign n_9701 =  n_9698 & ~n_9700;
assign n_9702 = ~n_9698 &  n_9700;
assign n_9703 = ~n_9701 & ~n_9702;
assign n_9704 =  x_2103 &  n_9703;
assign n_9705 = ~x_2103 & ~n_9703;
assign n_9706 =  n_8813 & ~n_9705;
assign n_9707 = ~n_9704 &  n_9706;
assign n_9708 =  x_1143 & ~n_8806;
assign n_9709 =  x_1623 & ~n_9662;
assign n_9710 = ~x_1623 &  n_9662;
assign n_9711 =  n_8824 & ~n_9710;
assign n_9712 = ~n_9709 &  n_9711;
assign n_9713 = ~n_9708 & ~n_9712;
assign n_9714 = ~n_9707 &  n_9713;
assign n_9715 = ~x_1815 &  n_9667;
assign n_9716 =  x_1815 & ~n_9667;
assign n_9717 = ~n_9715 & ~n_9716;
assign n_9718 = ~n_9671 & ~n_9675;
assign n_9719 =  n_9717 & ~n_9718;
assign n_9720 = ~n_9717 &  n_9718;
assign n_9721 = ~n_9719 & ~n_9720;
assign n_9722 = ~x_183 & ~n_9721;
assign n_9723 =  x_183 & ~n_9720;
assign n_9724 = ~n_9719 &  n_9723;
assign n_9725 =  n_8808 & ~n_9724;
assign n_9726 = ~n_9722 &  n_9725;
assign n_9727 = ~x_2007 &  n_9679;
assign n_9728 =  x_2007 & ~n_9679;
assign n_9729 = ~n_9727 & ~n_9728;
assign n_9730 = ~n_9683 & ~n_9687;
assign n_9731 =  n_9729 & ~n_9730;
assign n_9732 = ~n_9729 &  n_9730;
assign n_9733 = ~n_9731 & ~n_9732;
assign n_9734 = ~x_663 & ~n_9733;
assign n_9735 =  x_663 & ~n_9732;
assign n_9736 = ~n_9731 &  n_9735;
assign n_9737 =  n_8819 & ~n_9736;
assign n_9738 = ~n_9734 &  n_9737;
assign n_9739 = ~n_9726 & ~n_9738;
assign n_9740 =  n_9714 &  n_9739;
assign n_9741 =  x_1143 & ~n_9740;
assign n_9742 = ~x_1143 &  n_9740;
assign n_9743 = ~n_9741 & ~n_9742;
assign n_9744 = ~x_2774 &  n_9696;
assign n_9745 =  x_2774 & ~n_9696;
assign n_9746 = ~n_9744 & ~n_9745;
assign n_9747 =  x_2103 & ~n_9702;
assign n_9748 = ~n_9701 & ~n_9747;
assign n_9749 =  n_9746 & ~n_9748;
assign n_9750 = ~n_9746 &  n_9748;
assign n_9751 = ~n_9749 & ~n_9750;
assign n_9752 =  x_2102 &  n_9751;
assign n_9753 = ~x_2102 & ~n_9751;
assign n_9754 =  n_8813 & ~n_9753;
assign n_9755 = ~n_9752 &  n_9754;
assign n_9756 =  x_1142 & ~n_8806;
assign n_9757 =  x_1622 & ~n_9710;
assign n_9758 = ~x_1622 &  n_9710;
assign n_9759 =  n_8824 & ~n_9758;
assign n_9760 = ~n_9757 &  n_9759;
assign n_9761 = ~n_9756 & ~n_9760;
assign n_9762 = ~n_9755 &  n_9761;
assign n_9763 = ~x_1814 &  n_9715;
assign n_9764 =  x_1814 & ~n_9715;
assign n_9765 = ~n_9763 & ~n_9764;
assign n_9766 = ~n_9719 & ~n_9723;
assign n_9767 =  n_9765 & ~n_9766;
assign n_9768 = ~n_9765 &  n_9766;
assign n_9769 = ~n_9767 & ~n_9768;
assign n_9770 = ~x_182 & ~n_9769;
assign n_9771 =  x_182 & ~n_9768;
assign n_9772 = ~n_9767 &  n_9771;
assign n_9773 =  n_8808 & ~n_9772;
assign n_9774 = ~n_9770 &  n_9773;
assign n_9775 = ~x_2006 &  n_9727;
assign n_9776 =  x_2006 & ~n_9727;
assign n_9777 = ~n_9775 & ~n_9776;
assign n_9778 = ~n_9731 & ~n_9735;
assign n_9779 =  n_9777 & ~n_9778;
assign n_9780 = ~n_9777 &  n_9778;
assign n_9781 = ~n_9779 & ~n_9780;
assign n_9782 = ~x_662 & ~n_9781;
assign n_9783 =  x_662 & ~n_9780;
assign n_9784 = ~n_9779 &  n_9783;
assign n_9785 =  n_8819 & ~n_9784;
assign n_9786 = ~n_9782 &  n_9785;
assign n_9787 = ~n_9774 & ~n_9786;
assign n_9788 =  n_9762 &  n_9787;
assign n_9789 =  x_1142 & ~n_9788;
assign n_9790 = ~x_1142 &  n_9788;
assign n_9791 = ~n_9789 & ~n_9790;
assign n_9792 = ~x_2773 &  n_9744;
assign n_9793 =  x_2773 & ~n_9744;
assign n_9794 = ~n_9792 & ~n_9793;
assign n_9795 =  x_2102 & ~n_9750;
assign n_9796 = ~n_9749 & ~n_9795;
assign n_9797 =  n_9794 & ~n_9796;
assign n_9798 = ~n_9794 &  n_9796;
assign n_9799 = ~n_9797 & ~n_9798;
assign n_9800 =  x_2101 &  n_9799;
assign n_9801 = ~x_2101 & ~n_9799;
assign n_9802 =  n_8813 & ~n_9801;
assign n_9803 = ~n_9800 &  n_9802;
assign n_9804 =  x_1141 & ~n_8806;
assign n_9805 =  x_1621 & ~n_9758;
assign n_9806 = ~x_1621 &  n_9758;
assign n_9807 =  n_8824 & ~n_9806;
assign n_9808 = ~n_9805 &  n_9807;
assign n_9809 = ~n_9804 & ~n_9808;
assign n_9810 = ~n_9803 &  n_9809;
assign n_9811 = ~x_1813 &  n_9763;
assign n_9812 =  x_1813 & ~n_9763;
assign n_9813 = ~n_9811 & ~n_9812;
assign n_9814 = ~n_9767 & ~n_9771;
assign n_9815 =  n_9813 & ~n_9814;
assign n_9816 = ~n_9813 &  n_9814;
assign n_9817 = ~n_9815 & ~n_9816;
assign n_9818 = ~x_181 & ~n_9817;
assign n_9819 =  x_181 & ~n_9816;
assign n_9820 = ~n_9815 &  n_9819;
assign n_9821 =  n_8808 & ~n_9820;
assign n_9822 = ~n_9818 &  n_9821;
assign n_9823 = ~x_2005 &  n_9775;
assign n_9824 =  x_2005 & ~n_9775;
assign n_9825 = ~n_9823 & ~n_9824;
assign n_9826 = ~n_9779 & ~n_9783;
assign n_9827 =  n_9825 & ~n_9826;
assign n_9828 = ~n_9825 &  n_9826;
assign n_9829 = ~n_9827 & ~n_9828;
assign n_9830 = ~x_661 & ~n_9829;
assign n_9831 =  x_661 & ~n_9828;
assign n_9832 = ~n_9827 &  n_9831;
assign n_9833 =  n_8819 & ~n_9832;
assign n_9834 = ~n_9830 &  n_9833;
assign n_9835 = ~n_9822 & ~n_9834;
assign n_9836 =  n_9810 &  n_9835;
assign n_9837 =  x_1141 & ~n_9836;
assign n_9838 = ~x_1141 &  n_9836;
assign n_9839 = ~n_9837 & ~n_9838;
assign n_9840 = ~x_2772 &  n_9792;
assign n_9841 =  x_2772 & ~n_9792;
assign n_9842 = ~n_9840 & ~n_9841;
assign n_9843 =  x_2101 & ~n_9798;
assign n_9844 = ~n_9797 & ~n_9843;
assign n_9845 =  n_9842 & ~n_9844;
assign n_9846 = ~n_9842 &  n_9844;
assign n_9847 = ~n_9845 & ~n_9846;
assign n_9848 =  x_2100 &  n_9847;
assign n_9849 = ~x_2100 & ~n_9847;
assign n_9850 =  n_8813 & ~n_9849;
assign n_9851 = ~n_9848 &  n_9850;
assign n_9852 =  x_1140 & ~n_8806;
assign n_9853 =  x_1620 & ~n_9806;
assign n_9854 = ~x_1620 &  n_9806;
assign n_9855 =  n_8824 & ~n_9854;
assign n_9856 = ~n_9853 &  n_9855;
assign n_9857 = ~n_9852 & ~n_9856;
assign n_9858 = ~n_9851 &  n_9857;
assign n_9859 = ~x_1812 &  n_9811;
assign n_9860 =  x_1812 & ~n_9811;
assign n_9861 = ~n_9859 & ~n_9860;
assign n_9862 = ~n_9815 & ~n_9819;
assign n_9863 =  n_9861 & ~n_9862;
assign n_9864 = ~n_9861 &  n_9862;
assign n_9865 = ~n_9863 & ~n_9864;
assign n_9866 = ~x_180 & ~n_9865;
assign n_9867 =  x_180 & ~n_9864;
assign n_9868 = ~n_9863 &  n_9867;
assign n_9869 =  n_8808 & ~n_9868;
assign n_9870 = ~n_9866 &  n_9869;
assign n_9871 = ~x_2004 &  n_9823;
assign n_9872 =  x_2004 & ~n_9823;
assign n_9873 = ~n_9871 & ~n_9872;
assign n_9874 = ~n_9827 & ~n_9831;
assign n_9875 =  n_9873 & ~n_9874;
assign n_9876 = ~n_9873 &  n_9874;
assign n_9877 = ~n_9875 & ~n_9876;
assign n_9878 = ~x_660 & ~n_9877;
assign n_9879 =  x_660 & ~n_9876;
assign n_9880 = ~n_9875 &  n_9879;
assign n_9881 =  n_8819 & ~n_9880;
assign n_9882 = ~n_9878 &  n_9881;
assign n_9883 = ~n_9870 & ~n_9882;
assign n_9884 =  n_9858 &  n_9883;
assign n_9885 =  x_1140 & ~n_9884;
assign n_9886 = ~x_1140 &  n_9884;
assign n_9887 = ~n_9885 & ~n_9886;
assign n_9888 = ~x_2771 &  n_9840;
assign n_9889 =  x_2771 & ~n_9840;
assign n_9890 = ~n_9888 & ~n_9889;
assign n_9891 =  x_2100 & ~n_9846;
assign n_9892 = ~n_9845 & ~n_9891;
assign n_9893 =  n_9890 & ~n_9892;
assign n_9894 = ~n_9890 &  n_9892;
assign n_9895 = ~n_9893 & ~n_9894;
assign n_9896 =  x_2099 &  n_9895;
assign n_9897 = ~x_2099 & ~n_9895;
assign n_9898 =  n_8813 & ~n_9897;
assign n_9899 = ~n_9896 &  n_9898;
assign n_9900 =  x_1139 & ~n_8806;
assign n_9901 =  x_1619 & ~n_9854;
assign n_9902 = ~x_1619 &  n_9854;
assign n_9903 =  n_8824 & ~n_9902;
assign n_9904 = ~n_9901 &  n_9903;
assign n_9905 = ~n_9900 & ~n_9904;
assign n_9906 = ~n_9899 &  n_9905;
assign n_9907 = ~x_1811 &  n_9859;
assign n_9908 =  x_1811 & ~n_9859;
assign n_9909 = ~n_9907 & ~n_9908;
assign n_9910 = ~n_9863 & ~n_9867;
assign n_9911 =  n_9909 & ~n_9910;
assign n_9912 = ~n_9909 &  n_9910;
assign n_9913 = ~n_9911 & ~n_9912;
assign n_9914 = ~x_179 & ~n_9913;
assign n_9915 =  x_179 & ~n_9912;
assign n_9916 = ~n_9911 &  n_9915;
assign n_9917 =  n_8808 & ~n_9916;
assign n_9918 = ~n_9914 &  n_9917;
assign n_9919 = ~x_2003 &  n_9871;
assign n_9920 =  x_2003 & ~n_9871;
assign n_9921 = ~n_9919 & ~n_9920;
assign n_9922 = ~n_9875 & ~n_9879;
assign n_9923 =  n_9921 & ~n_9922;
assign n_9924 = ~n_9921 &  n_9922;
assign n_9925 = ~n_9923 & ~n_9924;
assign n_9926 = ~x_659 & ~n_9925;
assign n_9927 =  x_659 & ~n_9924;
assign n_9928 = ~n_9923 &  n_9927;
assign n_9929 =  n_8819 & ~n_9928;
assign n_9930 = ~n_9926 &  n_9929;
assign n_9931 = ~n_9918 & ~n_9930;
assign n_9932 =  n_9906 &  n_9931;
assign n_9933 =  x_1139 & ~n_9932;
assign n_9934 = ~x_1139 &  n_9932;
assign n_9935 = ~n_9933 & ~n_9934;
assign n_9936 = ~x_2770 &  n_9888;
assign n_9937 =  x_2770 & ~n_9888;
assign n_9938 = ~n_9936 & ~n_9937;
assign n_9939 =  x_2099 & ~n_9894;
assign n_9940 = ~n_9893 & ~n_9939;
assign n_9941 =  n_9938 & ~n_9940;
assign n_9942 = ~n_9938 &  n_9940;
assign n_9943 = ~n_9941 & ~n_9942;
assign n_9944 =  x_2098 &  n_9943;
assign n_9945 = ~x_2098 & ~n_9943;
assign n_9946 =  n_8813 & ~n_9945;
assign n_9947 = ~n_9944 &  n_9946;
assign n_9948 =  x_1138 & ~n_8806;
assign n_9949 =  x_1618 & ~n_9902;
assign n_9950 = ~x_1618 &  n_9902;
assign n_9951 =  n_8824 & ~n_9950;
assign n_9952 = ~n_9949 &  n_9951;
assign n_9953 = ~n_9948 & ~n_9952;
assign n_9954 = ~n_9947 &  n_9953;
assign n_9955 = ~x_1810 &  n_9907;
assign n_9956 =  x_1810 & ~n_9907;
assign n_9957 = ~n_9955 & ~n_9956;
assign n_9958 = ~n_9911 & ~n_9915;
assign n_9959 =  n_9957 & ~n_9958;
assign n_9960 = ~n_9957 &  n_9958;
assign n_9961 = ~n_9959 & ~n_9960;
assign n_9962 = ~x_178 & ~n_9961;
assign n_9963 =  x_178 & ~n_9960;
assign n_9964 = ~n_9959 &  n_9963;
assign n_9965 =  n_8808 & ~n_9964;
assign n_9966 = ~n_9962 &  n_9965;
assign n_9967 = ~x_2002 &  n_9919;
assign n_9968 =  x_2002 & ~n_9919;
assign n_9969 = ~n_9967 & ~n_9968;
assign n_9970 = ~n_9923 & ~n_9927;
assign n_9971 =  n_9969 & ~n_9970;
assign n_9972 = ~n_9969 &  n_9970;
assign n_9973 = ~n_9971 & ~n_9972;
assign n_9974 = ~x_658 & ~n_9973;
assign n_9975 =  x_658 & ~n_9972;
assign n_9976 = ~n_9971 &  n_9975;
assign n_9977 =  n_8819 & ~n_9976;
assign n_9978 = ~n_9974 &  n_9977;
assign n_9979 = ~n_9966 & ~n_9978;
assign n_9980 =  n_9954 &  n_9979;
assign n_9981 =  x_1138 & ~n_9980;
assign n_9982 = ~x_1138 &  n_9980;
assign n_9983 = ~n_9981 & ~n_9982;
assign n_9984 = ~x_2769 &  n_9936;
assign n_9985 =  x_2769 & ~n_9936;
assign n_9986 = ~n_9984 & ~n_9985;
assign n_9987 =  x_2098 & ~n_9942;
assign n_9988 = ~n_9941 & ~n_9987;
assign n_9989 =  n_9986 & ~n_9988;
assign n_9990 = ~n_9986 &  n_9988;
assign n_9991 = ~n_9989 & ~n_9990;
assign n_9992 =  x_2097 &  n_9991;
assign n_9993 = ~x_2097 & ~n_9991;
assign n_9994 =  n_8813 & ~n_9993;
assign n_9995 = ~n_9992 &  n_9994;
assign n_9996 =  x_1137 & ~n_8806;
assign n_9997 =  x_1617 & ~n_9950;
assign n_9998 = ~x_1617 &  n_9950;
assign n_9999 =  n_8824 & ~n_9998;
assign n_10000 = ~n_9997 &  n_9999;
assign n_10001 = ~n_9996 & ~n_10000;
assign n_10002 = ~n_9995 &  n_10001;
assign n_10003 = ~x_1809 &  n_9955;
assign n_10004 =  x_1809 & ~n_9955;
assign n_10005 = ~n_10003 & ~n_10004;
assign n_10006 = ~n_9959 & ~n_9963;
assign n_10007 =  n_10005 & ~n_10006;
assign n_10008 = ~n_10005 &  n_10006;
assign n_10009 = ~n_10007 & ~n_10008;
assign n_10010 = ~x_177 & ~n_10009;
assign n_10011 =  x_177 & ~n_10008;
assign n_10012 = ~n_10007 &  n_10011;
assign n_10013 =  n_8808 & ~n_10012;
assign n_10014 = ~n_10010 &  n_10013;
assign n_10015 = ~x_2001 &  n_9967;
assign n_10016 =  x_2001 & ~n_9967;
assign n_10017 = ~n_10015 & ~n_10016;
assign n_10018 = ~n_9971 & ~n_9975;
assign n_10019 =  n_10017 & ~n_10018;
assign n_10020 = ~n_10017 &  n_10018;
assign n_10021 = ~n_10019 & ~n_10020;
assign n_10022 = ~x_657 & ~n_10021;
assign n_10023 =  x_657 & ~n_10020;
assign n_10024 = ~n_10019 &  n_10023;
assign n_10025 =  n_8819 & ~n_10024;
assign n_10026 = ~n_10022 &  n_10025;
assign n_10027 = ~n_10014 & ~n_10026;
assign n_10028 =  n_10002 &  n_10027;
assign n_10029 =  x_1137 & ~n_10028;
assign n_10030 = ~x_1137 &  n_10028;
assign n_10031 = ~n_10029 & ~n_10030;
assign n_10032 = ~x_2768 &  n_9984;
assign n_10033 =  x_2768 & ~n_9984;
assign n_10034 = ~n_10032 & ~n_10033;
assign n_10035 =  x_2097 & ~n_9990;
assign n_10036 = ~n_9989 & ~n_10035;
assign n_10037 =  n_10034 & ~n_10036;
assign n_10038 = ~n_10034 &  n_10036;
assign n_10039 = ~n_10037 & ~n_10038;
assign n_10040 =  x_2096 &  n_10039;
assign n_10041 = ~x_2096 & ~n_10039;
assign n_10042 =  n_8813 & ~n_10041;
assign n_10043 = ~n_10040 &  n_10042;
assign n_10044 =  x_1136 & ~n_8806;
assign n_10045 =  x_1616 & ~n_9998;
assign n_10046 = ~x_1616 &  n_9998;
assign n_10047 =  n_8824 & ~n_10046;
assign n_10048 = ~n_10045 &  n_10047;
assign n_10049 = ~n_10044 & ~n_10048;
assign n_10050 = ~n_10043 &  n_10049;
assign n_10051 = ~x_1808 &  n_10003;
assign n_10052 =  x_1808 & ~n_10003;
assign n_10053 = ~n_10051 & ~n_10052;
assign n_10054 = ~n_10007 & ~n_10011;
assign n_10055 =  n_10053 & ~n_10054;
assign n_10056 = ~n_10053 &  n_10054;
assign n_10057 = ~n_10055 & ~n_10056;
assign n_10058 = ~x_176 & ~n_10057;
assign n_10059 =  x_176 & ~n_10056;
assign n_10060 = ~n_10055 &  n_10059;
assign n_10061 =  n_8808 & ~n_10060;
assign n_10062 = ~n_10058 &  n_10061;
assign n_10063 = ~x_2000 &  n_10015;
assign n_10064 =  x_2000 & ~n_10015;
assign n_10065 = ~n_10063 & ~n_10064;
assign n_10066 = ~n_10019 & ~n_10023;
assign n_10067 =  n_10065 & ~n_10066;
assign n_10068 = ~n_10065 &  n_10066;
assign n_10069 = ~n_10067 & ~n_10068;
assign n_10070 = ~x_656 & ~n_10069;
assign n_10071 =  x_656 & ~n_10068;
assign n_10072 = ~n_10067 &  n_10071;
assign n_10073 =  n_8819 & ~n_10072;
assign n_10074 = ~n_10070 &  n_10073;
assign n_10075 = ~n_10062 & ~n_10074;
assign n_10076 =  n_10050 &  n_10075;
assign n_10077 =  x_1136 & ~n_10076;
assign n_10078 = ~x_1136 &  n_10076;
assign n_10079 = ~n_10077 & ~n_10078;
assign n_10080 = ~x_2767 &  n_10032;
assign n_10081 =  x_2767 & ~n_10032;
assign n_10082 = ~n_10080 & ~n_10081;
assign n_10083 =  x_2096 & ~n_10038;
assign n_10084 = ~n_10037 & ~n_10083;
assign n_10085 =  n_10082 & ~n_10084;
assign n_10086 = ~n_10082 &  n_10084;
assign n_10087 = ~n_10085 & ~n_10086;
assign n_10088 =  x_2095 &  n_10087;
assign n_10089 = ~x_2095 & ~n_10087;
assign n_10090 =  n_8813 & ~n_10089;
assign n_10091 = ~n_10088 &  n_10090;
assign n_10092 =  x_1135 & ~n_8806;
assign n_10093 =  x_1615 & ~n_10046;
assign n_10094 = ~x_1615 &  n_10046;
assign n_10095 =  n_8824 & ~n_10094;
assign n_10096 = ~n_10093 &  n_10095;
assign n_10097 = ~n_10092 & ~n_10096;
assign n_10098 = ~n_10091 &  n_10097;
assign n_10099 = ~x_1807 &  n_10051;
assign n_10100 =  x_1807 & ~n_10051;
assign n_10101 = ~n_10099 & ~n_10100;
assign n_10102 = ~n_10055 & ~n_10059;
assign n_10103 =  n_10101 & ~n_10102;
assign n_10104 = ~n_10101 &  n_10102;
assign n_10105 = ~n_10103 & ~n_10104;
assign n_10106 = ~x_175 & ~n_10105;
assign n_10107 =  x_175 & ~n_10104;
assign n_10108 = ~n_10103 &  n_10107;
assign n_10109 =  n_8808 & ~n_10108;
assign n_10110 = ~n_10106 &  n_10109;
assign n_10111 = ~x_1999 &  n_10063;
assign n_10112 =  x_1999 & ~n_10063;
assign n_10113 = ~n_10111 & ~n_10112;
assign n_10114 = ~n_10067 & ~n_10071;
assign n_10115 =  n_10113 & ~n_10114;
assign n_10116 = ~n_10113 &  n_10114;
assign n_10117 = ~n_10115 & ~n_10116;
assign n_10118 = ~x_655 & ~n_10117;
assign n_10119 =  x_655 & ~n_10116;
assign n_10120 = ~n_10115 &  n_10119;
assign n_10121 =  n_8819 & ~n_10120;
assign n_10122 = ~n_10118 &  n_10121;
assign n_10123 = ~n_10110 & ~n_10122;
assign n_10124 =  n_10098 &  n_10123;
assign n_10125 =  x_1135 & ~n_10124;
assign n_10126 = ~x_1135 &  n_10124;
assign n_10127 = ~n_10125 & ~n_10126;
assign n_10128 = ~x_2766 &  n_10080;
assign n_10129 =  x_2766 & ~n_10080;
assign n_10130 = ~n_10128 & ~n_10129;
assign n_10131 =  x_2095 & ~n_10086;
assign n_10132 = ~n_10085 & ~n_10131;
assign n_10133 =  n_10130 & ~n_10132;
assign n_10134 = ~n_10130 &  n_10132;
assign n_10135 = ~n_10133 & ~n_10134;
assign n_10136 =  x_2094 &  n_10135;
assign n_10137 = ~x_2094 & ~n_10135;
assign n_10138 =  n_8813 & ~n_10137;
assign n_10139 = ~n_10136 &  n_10138;
assign n_10140 =  x_1134 & ~n_8806;
assign n_10141 =  x_1614 & ~n_10094;
assign n_10142 = ~x_1614 &  n_10094;
assign n_10143 =  n_8824 & ~n_10142;
assign n_10144 = ~n_10141 &  n_10143;
assign n_10145 = ~n_10140 & ~n_10144;
assign n_10146 = ~n_10139 &  n_10145;
assign n_10147 = ~x_1806 &  n_10099;
assign n_10148 =  x_1806 & ~n_10099;
assign n_10149 = ~n_10147 & ~n_10148;
assign n_10150 = ~n_10103 & ~n_10107;
assign n_10151 =  n_10149 & ~n_10150;
assign n_10152 = ~n_10149 &  n_10150;
assign n_10153 = ~n_10151 & ~n_10152;
assign n_10154 = ~x_174 & ~n_10153;
assign n_10155 =  x_174 & ~n_10152;
assign n_10156 = ~n_10151 &  n_10155;
assign n_10157 =  n_8808 & ~n_10156;
assign n_10158 = ~n_10154 &  n_10157;
assign n_10159 = ~x_1998 &  n_10111;
assign n_10160 =  x_1998 & ~n_10111;
assign n_10161 = ~n_10159 & ~n_10160;
assign n_10162 = ~n_10115 & ~n_10119;
assign n_10163 =  n_10161 & ~n_10162;
assign n_10164 = ~n_10161 &  n_10162;
assign n_10165 = ~n_10163 & ~n_10164;
assign n_10166 = ~x_654 & ~n_10165;
assign n_10167 =  x_654 & ~n_10164;
assign n_10168 = ~n_10163 &  n_10167;
assign n_10169 =  n_8819 & ~n_10168;
assign n_10170 = ~n_10166 &  n_10169;
assign n_10171 = ~n_10158 & ~n_10170;
assign n_10172 =  n_10146 &  n_10171;
assign n_10173 =  x_1134 & ~n_10172;
assign n_10174 = ~x_1134 &  n_10172;
assign n_10175 = ~n_10173 & ~n_10174;
assign n_10176 = ~x_2765 &  n_10128;
assign n_10177 =  x_2765 & ~n_10128;
assign n_10178 = ~n_10176 & ~n_10177;
assign n_10179 =  x_2094 & ~n_10134;
assign n_10180 = ~n_10133 & ~n_10179;
assign n_10181 =  n_10178 & ~n_10180;
assign n_10182 = ~n_10178 &  n_10180;
assign n_10183 = ~n_10181 & ~n_10182;
assign n_10184 =  x_2093 &  n_10183;
assign n_10185 = ~x_2093 & ~n_10183;
assign n_10186 =  n_8813 & ~n_10185;
assign n_10187 = ~n_10184 &  n_10186;
assign n_10188 =  x_1133 & ~n_8806;
assign n_10189 =  x_1613 & ~n_10142;
assign n_10190 = ~x_1613 &  n_10142;
assign n_10191 =  n_8824 & ~n_10190;
assign n_10192 = ~n_10189 &  n_10191;
assign n_10193 = ~n_10188 & ~n_10192;
assign n_10194 = ~n_10187 &  n_10193;
assign n_10195 = ~x_1805 &  n_10147;
assign n_10196 =  x_1805 & ~n_10147;
assign n_10197 = ~n_10195 & ~n_10196;
assign n_10198 = ~n_10151 & ~n_10155;
assign n_10199 =  n_10197 & ~n_10198;
assign n_10200 = ~n_10197 &  n_10198;
assign n_10201 = ~n_10199 & ~n_10200;
assign n_10202 = ~x_173 & ~n_10201;
assign n_10203 =  x_173 & ~n_10200;
assign n_10204 = ~n_10199 &  n_10203;
assign n_10205 =  n_8808 & ~n_10204;
assign n_10206 = ~n_10202 &  n_10205;
assign n_10207 = ~x_1997 &  n_10159;
assign n_10208 =  x_1997 & ~n_10159;
assign n_10209 = ~n_10207 & ~n_10208;
assign n_10210 = ~n_10163 & ~n_10167;
assign n_10211 =  n_10209 & ~n_10210;
assign n_10212 = ~n_10209 &  n_10210;
assign n_10213 = ~n_10211 & ~n_10212;
assign n_10214 = ~x_653 & ~n_10213;
assign n_10215 =  x_653 & ~n_10212;
assign n_10216 = ~n_10211 &  n_10215;
assign n_10217 =  n_8819 & ~n_10216;
assign n_10218 = ~n_10214 &  n_10217;
assign n_10219 = ~n_10206 & ~n_10218;
assign n_10220 =  n_10194 &  n_10219;
assign n_10221 =  x_1133 & ~n_10220;
assign n_10222 = ~x_1133 &  n_10220;
assign n_10223 = ~n_10221 & ~n_10222;
assign n_10224 = ~x_2764 &  n_10176;
assign n_10225 =  x_2764 & ~n_10176;
assign n_10226 = ~n_10224 & ~n_10225;
assign n_10227 =  x_2093 & ~n_10182;
assign n_10228 = ~n_10181 & ~n_10227;
assign n_10229 =  n_10226 & ~n_10228;
assign n_10230 = ~n_10226 &  n_10228;
assign n_10231 = ~n_10229 & ~n_10230;
assign n_10232 =  x_2092 &  n_10231;
assign n_10233 = ~x_2092 & ~n_10231;
assign n_10234 =  n_8813 & ~n_10233;
assign n_10235 = ~n_10232 &  n_10234;
assign n_10236 =  x_1132 & ~n_8806;
assign n_10237 =  x_1612 & ~n_10190;
assign n_10238 = ~x_1612 &  n_10190;
assign n_10239 =  n_8824 & ~n_10238;
assign n_10240 = ~n_10237 &  n_10239;
assign n_10241 = ~n_10236 & ~n_10240;
assign n_10242 = ~n_10235 &  n_10241;
assign n_10243 = ~x_1804 &  n_10195;
assign n_10244 =  x_1804 & ~n_10195;
assign n_10245 = ~n_10243 & ~n_10244;
assign n_10246 = ~n_10199 & ~n_10203;
assign n_10247 =  n_10245 & ~n_10246;
assign n_10248 = ~n_10245 &  n_10246;
assign n_10249 = ~n_10247 & ~n_10248;
assign n_10250 = ~x_172 & ~n_10249;
assign n_10251 =  x_172 & ~n_10248;
assign n_10252 = ~n_10247 &  n_10251;
assign n_10253 =  n_8808 & ~n_10252;
assign n_10254 = ~n_10250 &  n_10253;
assign n_10255 = ~x_1996 &  n_10207;
assign n_10256 =  x_1996 & ~n_10207;
assign n_10257 = ~n_10255 & ~n_10256;
assign n_10258 = ~n_10211 & ~n_10215;
assign n_10259 =  n_10257 & ~n_10258;
assign n_10260 = ~n_10257 &  n_10258;
assign n_10261 = ~n_10259 & ~n_10260;
assign n_10262 = ~x_652 & ~n_10261;
assign n_10263 =  x_652 & ~n_10260;
assign n_10264 = ~n_10259 &  n_10263;
assign n_10265 =  n_8819 & ~n_10264;
assign n_10266 = ~n_10262 &  n_10265;
assign n_10267 = ~n_10254 & ~n_10266;
assign n_10268 =  n_10242 &  n_10267;
assign n_10269 =  x_1132 & ~n_10268;
assign n_10270 = ~x_1132 &  n_10268;
assign n_10271 = ~n_10269 & ~n_10270;
assign n_10272 = ~n_10247 & ~n_10251;
assign n_10273 =  x_171 & ~x_1803;
assign n_10274 = ~x_171 &  x_1803;
assign n_10275 = ~n_10273 & ~n_10274;
assign n_10276 =  n_10243 &  n_10275;
assign n_10277 = ~n_10243 & ~n_10275;
assign n_10278 = ~n_10276 & ~n_10277;
assign n_10279 =  n_10272 & ~n_10278;
assign n_10280 = ~n_10272 &  n_10278;
assign n_10281 =  n_8808 & ~n_10280;
assign n_10282 = ~n_10279 &  n_10281;
assign n_10283 =  x_1131 & ~n_8806;
assign n_10284 = ~x_1611 &  n_10238;
assign n_10285 =  x_1611 & ~n_10238;
assign n_10286 =  n_8824 & ~n_10285;
assign n_10287 = ~n_10284 &  n_10286;
assign n_10288 = ~n_10283 & ~n_10287;
assign n_10289 = ~n_10282 &  n_10288;
assign n_10290 = ~n_10259 & ~n_10263;
assign n_10291 =  x_651 & ~x_1995;
assign n_10292 = ~x_651 &  x_1995;
assign n_10293 = ~n_10291 & ~n_10292;
assign n_10294 =  n_10255 &  n_10293;
assign n_10295 = ~n_10255 & ~n_10293;
assign n_10296 = ~n_10294 & ~n_10295;
assign n_10297 =  n_10290 & ~n_10296;
assign n_10298 = ~n_10290 &  n_10296;
assign n_10299 =  n_8819 & ~n_10298;
assign n_10300 = ~n_10297 &  n_10299;
assign n_10301 =  x_2092 & ~n_10230;
assign n_10302 = ~n_10229 & ~n_10301;
assign n_10303 =  x_2091 & ~x_2763;
assign n_10304 = ~x_2091 &  x_2763;
assign n_10305 = ~n_10303 & ~n_10304;
assign n_10306 =  n_10224 &  n_10305;
assign n_10307 = ~n_10224 & ~n_10305;
assign n_10308 = ~n_10306 & ~n_10307;
assign n_10309 =  n_10302 & ~n_10308;
assign n_10310 = ~n_10302 &  n_10308;
assign n_10311 =  n_8813 & ~n_10310;
assign n_10312 = ~n_10309 &  n_10311;
assign n_10313 = ~n_10300 & ~n_10312;
assign n_10314 =  n_10289 &  n_10313;
assign n_10315 =  x_1131 & ~n_10314;
assign n_10316 = ~x_1131 &  n_10314;
assign n_10317 = ~n_10315 & ~n_10316;
assign n_10318 =  x_42 &  n_1314;
assign n_10319 =  x_39 &  n_187;
assign n_10320 =  n_10319 &  n_982;
assign n_10321 = ~n_10320 & ~n_3862;
assign n_10322 =  n_10318 & ~n_10321;
assign n_10323 =  x_1130 & ~n_10322;
assign n_10324 =  i_32 &  n_10322;
assign n_10325 = ~n_10323 & ~n_10324;
assign n_10326 =  x_1130 & ~n_10325;
assign n_10327 = ~x_1130 &  n_10325;
assign n_10328 = ~n_10326 & ~n_10327;
assign n_10329 =  x_1129 & ~n_10322;
assign n_10330 =  i_31 &  n_10322;
assign n_10331 = ~n_10329 & ~n_10330;
assign n_10332 =  x_1129 & ~n_10331;
assign n_10333 = ~x_1129 &  n_10331;
assign n_10334 = ~n_10332 & ~n_10333;
assign n_10335 =  x_1128 & ~n_10322;
assign n_10336 =  i_30 &  n_10322;
assign n_10337 = ~n_10335 & ~n_10336;
assign n_10338 =  x_1128 & ~n_10337;
assign n_10339 = ~x_1128 &  n_10337;
assign n_10340 = ~n_10338 & ~n_10339;
assign n_10341 =  x_1127 & ~n_10322;
assign n_10342 =  i_29 &  n_10322;
assign n_10343 = ~n_10341 & ~n_10342;
assign n_10344 =  x_1127 & ~n_10343;
assign n_10345 = ~x_1127 &  n_10343;
assign n_10346 = ~n_10344 & ~n_10345;
assign n_10347 =  x_1126 & ~n_10322;
assign n_10348 =  i_28 &  n_10322;
assign n_10349 = ~n_10347 & ~n_10348;
assign n_10350 =  x_1126 & ~n_10349;
assign n_10351 = ~x_1126 &  n_10349;
assign n_10352 = ~n_10350 & ~n_10351;
assign n_10353 =  x_1125 & ~n_10322;
assign n_10354 =  i_27 &  n_10322;
assign n_10355 = ~n_10353 & ~n_10354;
assign n_10356 =  x_1125 & ~n_10355;
assign n_10357 = ~x_1125 &  n_10355;
assign n_10358 = ~n_10356 & ~n_10357;
assign n_10359 =  x_1124 & ~n_10322;
assign n_10360 =  i_26 &  n_10322;
assign n_10361 = ~n_10359 & ~n_10360;
assign n_10362 =  x_1124 & ~n_10361;
assign n_10363 = ~x_1124 &  n_10361;
assign n_10364 = ~n_10362 & ~n_10363;
assign n_10365 =  x_1123 & ~n_10322;
assign n_10366 =  i_25 &  n_10322;
assign n_10367 = ~n_10365 & ~n_10366;
assign n_10368 =  x_1123 & ~n_10367;
assign n_10369 = ~x_1123 &  n_10367;
assign n_10370 = ~n_10368 & ~n_10369;
assign n_10371 =  x_1122 & ~n_10322;
assign n_10372 =  i_24 &  n_10322;
assign n_10373 = ~n_10371 & ~n_10372;
assign n_10374 =  x_1122 & ~n_10373;
assign n_10375 = ~x_1122 &  n_10373;
assign n_10376 = ~n_10374 & ~n_10375;
assign n_10377 =  x_1121 & ~n_10322;
assign n_10378 =  i_23 &  n_10322;
assign n_10379 = ~n_10377 & ~n_10378;
assign n_10380 =  x_1121 & ~n_10379;
assign n_10381 = ~x_1121 &  n_10379;
assign n_10382 = ~n_10380 & ~n_10381;
assign n_10383 =  x_1120 & ~n_10322;
assign n_10384 =  i_22 &  n_10322;
assign n_10385 = ~n_10383 & ~n_10384;
assign n_10386 =  x_1120 & ~n_10385;
assign n_10387 = ~x_1120 &  n_10385;
assign n_10388 = ~n_10386 & ~n_10387;
assign n_10389 =  x_1119 & ~n_10322;
assign n_10390 =  i_21 &  n_10322;
assign n_10391 = ~n_10389 & ~n_10390;
assign n_10392 =  x_1119 & ~n_10391;
assign n_10393 = ~x_1119 &  n_10391;
assign n_10394 = ~n_10392 & ~n_10393;
assign n_10395 =  x_1118 & ~n_10322;
assign n_10396 =  i_20 &  n_10322;
assign n_10397 = ~n_10395 & ~n_10396;
assign n_10398 =  x_1118 & ~n_10397;
assign n_10399 = ~x_1118 &  n_10397;
assign n_10400 = ~n_10398 & ~n_10399;
assign n_10401 =  x_1117 & ~n_10322;
assign n_10402 =  i_19 &  n_10322;
assign n_10403 = ~n_10401 & ~n_10402;
assign n_10404 =  x_1117 & ~n_10403;
assign n_10405 = ~x_1117 &  n_10403;
assign n_10406 = ~n_10404 & ~n_10405;
assign n_10407 =  x_1116 & ~n_10322;
assign n_10408 =  i_18 &  n_10322;
assign n_10409 = ~n_10407 & ~n_10408;
assign n_10410 =  x_1116 & ~n_10409;
assign n_10411 = ~x_1116 &  n_10409;
assign n_10412 = ~n_10410 & ~n_10411;
assign n_10413 =  x_1115 & ~n_10322;
assign n_10414 =  i_17 &  n_10322;
assign n_10415 = ~n_10413 & ~n_10414;
assign n_10416 =  x_1115 & ~n_10415;
assign n_10417 = ~x_1115 &  n_10415;
assign n_10418 = ~n_10416 & ~n_10417;
assign n_10419 =  x_1114 & ~n_10322;
assign n_10420 =  i_16 &  n_10322;
assign n_10421 = ~n_10419 & ~n_10420;
assign n_10422 =  x_1114 & ~n_10421;
assign n_10423 = ~x_1114 &  n_10421;
assign n_10424 = ~n_10422 & ~n_10423;
assign n_10425 =  x_1113 & ~n_10322;
assign n_10426 =  i_15 &  n_10322;
assign n_10427 = ~n_10425 & ~n_10426;
assign n_10428 =  x_1113 & ~n_10427;
assign n_10429 = ~x_1113 &  n_10427;
assign n_10430 = ~n_10428 & ~n_10429;
assign n_10431 =  x_1112 & ~n_10322;
assign n_10432 =  i_14 &  n_10322;
assign n_10433 = ~n_10431 & ~n_10432;
assign n_10434 =  x_1112 & ~n_10433;
assign n_10435 = ~x_1112 &  n_10433;
assign n_10436 = ~n_10434 & ~n_10435;
assign n_10437 =  x_1111 & ~n_10322;
assign n_10438 =  i_13 &  n_10322;
assign n_10439 = ~n_10437 & ~n_10438;
assign n_10440 =  x_1111 & ~n_10439;
assign n_10441 = ~x_1111 &  n_10439;
assign n_10442 = ~n_10440 & ~n_10441;
assign n_10443 =  x_1110 & ~n_10322;
assign n_10444 =  i_12 &  n_10322;
assign n_10445 = ~n_10443 & ~n_10444;
assign n_10446 =  x_1110 & ~n_10445;
assign n_10447 = ~x_1110 &  n_10445;
assign n_10448 = ~n_10446 & ~n_10447;
assign n_10449 =  x_1109 & ~n_10322;
assign n_10450 =  i_11 &  n_10322;
assign n_10451 = ~n_10449 & ~n_10450;
assign n_10452 =  x_1109 & ~n_10451;
assign n_10453 = ~x_1109 &  n_10451;
assign n_10454 = ~n_10452 & ~n_10453;
assign n_10455 =  x_1108 & ~n_10322;
assign n_10456 =  i_10 &  n_10322;
assign n_10457 = ~n_10455 & ~n_10456;
assign n_10458 =  x_1108 & ~n_10457;
assign n_10459 = ~x_1108 &  n_10457;
assign n_10460 = ~n_10458 & ~n_10459;
assign n_10461 =  x_1107 & ~n_10322;
assign n_10462 =  i_9 &  n_10322;
assign n_10463 = ~n_10461 & ~n_10462;
assign n_10464 =  x_1107 & ~n_10463;
assign n_10465 = ~x_1107 &  n_10463;
assign n_10466 = ~n_10464 & ~n_10465;
assign n_10467 =  x_1106 & ~n_10322;
assign n_10468 =  i_8 &  n_10322;
assign n_10469 = ~n_10467 & ~n_10468;
assign n_10470 =  x_1106 & ~n_10469;
assign n_10471 = ~x_1106 &  n_10469;
assign n_10472 = ~n_10470 & ~n_10471;
assign n_10473 =  x_1105 & ~n_10322;
assign n_10474 =  i_7 &  n_10322;
assign n_10475 = ~n_10473 & ~n_10474;
assign n_10476 =  x_1105 & ~n_10475;
assign n_10477 = ~x_1105 &  n_10475;
assign n_10478 = ~n_10476 & ~n_10477;
assign n_10479 =  x_1104 & ~n_10322;
assign n_10480 =  i_6 &  n_10322;
assign n_10481 = ~n_10479 & ~n_10480;
assign n_10482 =  x_1104 & ~n_10481;
assign n_10483 = ~x_1104 &  n_10481;
assign n_10484 = ~n_10482 & ~n_10483;
assign n_10485 =  x_1103 & ~n_10322;
assign n_10486 =  i_5 &  n_10322;
assign n_10487 = ~n_10485 & ~n_10486;
assign n_10488 =  x_1103 & ~n_10487;
assign n_10489 = ~x_1103 &  n_10487;
assign n_10490 = ~n_10488 & ~n_10489;
assign n_10491 =  x_1102 & ~n_10322;
assign n_10492 =  i_4 &  n_10322;
assign n_10493 = ~n_10491 & ~n_10492;
assign n_10494 =  x_1102 & ~n_10493;
assign n_10495 = ~x_1102 &  n_10493;
assign n_10496 = ~n_10494 & ~n_10495;
assign n_10497 =  x_1101 & ~n_10322;
assign n_10498 =  i_3 &  n_10322;
assign n_10499 = ~n_10497 & ~n_10498;
assign n_10500 =  x_1101 & ~n_10499;
assign n_10501 = ~x_1101 &  n_10499;
assign n_10502 = ~n_10500 & ~n_10501;
assign n_10503 =  x_1100 & ~n_10322;
assign n_10504 =  i_2 &  n_10322;
assign n_10505 = ~n_10503 & ~n_10504;
assign n_10506 =  x_1100 & ~n_10505;
assign n_10507 = ~x_1100 &  n_10505;
assign n_10508 = ~n_10506 & ~n_10507;
assign n_10509 =  x_1099 & ~n_10322;
assign n_10510 =  i_1 &  n_10322;
assign n_10511 = ~n_10509 & ~n_10510;
assign n_10512 =  x_1099 & ~n_10511;
assign n_10513 = ~x_1099 &  n_10511;
assign n_10514 = ~n_10512 & ~n_10513;
assign n_10515 =  x_39 &  n_3275;
assign n_10516 =  n_1706 &  n_10515;
assign n_10517 =  x_40 &  n_10516;
assign n_10518 =  n_10319 &  n_190;
assign n_10519 =  n_3858 &  n_10518;
assign n_10520 = ~n_10517 & ~n_10519;
assign n_10521 =  n_184 &  n_4057;
assign n_10522 =  n_4992 &  n_10521;
assign n_10523 =  n_8818 &  n_191;
assign n_10524 = ~n_10522 & ~n_10523;
assign n_10525 =  n_10520 &  n_10524;
assign n_10526 =  x_1098 &  n_10525;
assign n_10527 =  x_874 &  n_10517;
assign n_10528 =  x_266 &  x_1706;
assign n_10529 = ~x_266 & ~x_1706;
assign n_10530 = ~n_10528 & ~n_10529;
assign n_10531 =  n_10522 &  n_10530;
assign n_10532 =  x_458 &  x_2346;
assign n_10533 = ~x_458 & ~x_2346;
assign n_10534 = ~n_10532 & ~n_10533;
assign n_10535 =  n_10523 &  n_10534;
assign n_10536 =  x_234 &  x_2698;
assign n_10537 = ~x_234 & ~x_2698;
assign n_10538 = ~n_10536 & ~n_10537;
assign n_10539 =  n_10519 &  n_10538;
assign n_10540 = ~n_10535 & ~n_10539;
assign n_10541 = ~n_10531 &  n_10540;
assign n_10542 = ~n_10527 &  n_10541;
assign n_10543 = ~n_10526 &  n_10542;
assign n_10544 =  x_1098 & ~n_10543;
assign n_10545 = ~x_1098 &  n_10543;
assign n_10546 = ~n_10544 & ~n_10545;
assign n_10547 =  x_1097 &  n_10525;
assign n_10548 = ~x_233 & ~x_234;
assign n_10549 =  x_233 &  x_234;
assign n_10550 = ~n_10548 & ~n_10549;
assign n_10551 =  x_2697 &  n_10550;
assign n_10552 = ~x_2697 & ~n_10550;
assign n_10553 = ~n_10551 & ~n_10552;
assign n_10554 = ~n_10536 & ~n_10553;
assign n_10555 =  n_10536 &  n_10553;
assign n_10556 =  n_10519 & ~n_10555;
assign n_10557 = ~n_10554 &  n_10556;
assign n_10558 = ~x_1705 & ~x_1706;
assign n_10559 =  x_1705 &  x_1706;
assign n_10560 = ~n_10558 & ~n_10559;
assign n_10561 =  x_265 &  n_10560;
assign n_10562 = ~x_265 & ~n_10560;
assign n_10563 = ~n_10561 & ~n_10562;
assign n_10564 = ~n_10528 & ~n_10563;
assign n_10565 =  n_10528 &  n_10563;
assign n_10566 =  n_10522 & ~n_10565;
assign n_10567 = ~n_10564 &  n_10566;
assign n_10568 = ~n_10557 & ~n_10567;
assign n_10569 = ~x_2345 & ~x_2346;
assign n_10570 =  x_2345 &  x_2346;
assign n_10571 = ~n_10569 & ~n_10570;
assign n_10572 =  x_457 &  n_10571;
assign n_10573 = ~x_457 & ~n_10571;
assign n_10574 = ~n_10572 & ~n_10573;
assign n_10575 = ~n_10532 & ~n_10574;
assign n_10576 =  n_10532 &  n_10574;
assign n_10577 =  n_10523 & ~n_10576;
assign n_10578 = ~n_10575 &  n_10577;
assign n_10579 = ~x_873 & ~x_874;
assign n_10580 =  x_873 &  x_874;
assign n_10581 = ~n_10579 & ~n_10580;
assign n_10582 =  n_10517 &  n_10581;
assign n_10583 = ~n_10578 & ~n_10582;
assign n_10584 =  n_10568 &  n_10583;
assign n_10585 = ~n_10547 &  n_10584;
assign n_10586 =  x_1097 & ~n_10585;
assign n_10587 = ~x_1097 &  n_10585;
assign n_10588 = ~n_10586 & ~n_10587;
assign n_10589 = ~x_2344 &  n_10569;
assign n_10590 =  x_2344 & ~n_10569;
assign n_10591 = ~n_10589 & ~n_10590;
assign n_10592 = ~x_457 &  x_2345;
assign n_10593 =  n_10532 & ~n_10592;
assign n_10594 = ~n_10593 & ~n_10572;
assign n_10595 =  n_10591 & ~n_10594;
assign n_10596 = ~n_10591 &  n_10594;
assign n_10597 = ~n_10595 & ~n_10596;
assign n_10598 = ~x_456 & ~n_10597;
assign n_10599 =  x_456 & ~n_10596;
assign n_10600 = ~n_10595 &  n_10599;
assign n_10601 =  n_10523 & ~n_10600;
assign n_10602 = ~n_10598 &  n_10601;
assign n_10603 = ~x_872 &  n_10579;
assign n_10604 =  x_872 & ~n_10579;
assign n_10605 = ~n_10603 & ~n_10604;
assign n_10606 =  n_10517 &  n_10605;
assign n_10607 = ~n_10602 & ~n_10606;
assign n_10608 = ~x_1704 &  n_10558;
assign n_10609 =  x_1704 & ~n_10558;
assign n_10610 = ~n_10608 & ~n_10609;
assign n_10611 = ~x_265 &  x_1705;
assign n_10612 =  n_10528 & ~n_10611;
assign n_10613 = ~n_10612 & ~n_10561;
assign n_10614 =  n_10610 & ~n_10613;
assign n_10615 = ~n_10610 &  n_10613;
assign n_10616 = ~n_10614 & ~n_10615;
assign n_10617 = ~x_264 & ~n_10616;
assign n_10618 =  x_264 & ~n_10615;
assign n_10619 = ~n_10614 &  n_10618;
assign n_10620 =  n_10522 & ~n_10619;
assign n_10621 = ~n_10617 &  n_10620;
assign n_10622 = ~x_232 &  n_10548;
assign n_10623 =  x_232 & ~n_10548;
assign n_10624 = ~n_10622 & ~n_10623;
assign n_10625 =  x_233 & ~x_2697;
assign n_10626 =  n_10536 & ~n_10625;
assign n_10627 = ~n_10626 & ~n_10551;
assign n_10628 =  n_10624 & ~n_10627;
assign n_10629 = ~n_10624 &  n_10627;
assign n_10630 = ~n_10628 & ~n_10629;
assign n_10631 = ~x_2696 & ~n_10630;
assign n_10632 =  x_2696 & ~n_10629;
assign n_10633 = ~n_10628 &  n_10632;
assign n_10634 =  n_10519 & ~n_10633;
assign n_10635 = ~n_10631 &  n_10634;
assign n_10636 =  x_1096 &  n_10525;
assign n_10637 = ~n_10635 & ~n_10636;
assign n_10638 = ~n_10621 &  n_10637;
assign n_10639 =  n_10607 &  n_10638;
assign n_10640 =  x_1096 & ~n_10639;
assign n_10641 = ~x_1096 &  n_10639;
assign n_10642 = ~n_10640 & ~n_10641;
assign n_10643 = ~x_231 &  n_10622;
assign n_10644 =  x_231 & ~n_10622;
assign n_10645 = ~n_10643 & ~n_10644;
assign n_10646 = ~n_10628 & ~n_10632;
assign n_10647 =  n_10645 & ~n_10646;
assign n_10648 = ~n_10645 &  n_10646;
assign n_10649 = ~n_10647 & ~n_10648;
assign n_10650 = ~x_2695 & ~n_10649;
assign n_10651 =  x_2695 & ~n_10648;
assign n_10652 = ~n_10647 &  n_10651;
assign n_10653 =  n_10519 & ~n_10652;
assign n_10654 = ~n_10650 &  n_10653;
assign n_10655 =  x_1095 &  n_10525;
assign n_10656 = ~x_871 &  n_10603;
assign n_10657 =  x_871 & ~n_10603;
assign n_10658 = ~n_10656 & ~n_10657;
assign n_10659 =  n_10517 &  n_10658;
assign n_10660 = ~n_10655 & ~n_10659;
assign n_10661 = ~n_10654 &  n_10660;
assign n_10662 = ~x_2343 &  n_10589;
assign n_10663 =  x_2343 & ~n_10589;
assign n_10664 = ~n_10662 & ~n_10663;
assign n_10665 = ~n_10595 & ~n_10599;
assign n_10666 =  n_10664 & ~n_10665;
assign n_10667 = ~n_10664 &  n_10665;
assign n_10668 = ~n_10666 & ~n_10667;
assign n_10669 = ~x_455 & ~n_10668;
assign n_10670 =  x_455 & ~n_10667;
assign n_10671 = ~n_10666 &  n_10670;
assign n_10672 =  n_10523 & ~n_10671;
assign n_10673 = ~n_10669 &  n_10672;
assign n_10674 = ~x_1703 &  n_10608;
assign n_10675 =  x_1703 & ~n_10608;
assign n_10676 = ~n_10674 & ~n_10675;
assign n_10677 = ~n_10614 & ~n_10618;
assign n_10678 =  n_10676 & ~n_10677;
assign n_10679 = ~n_10676 &  n_10677;
assign n_10680 = ~n_10678 & ~n_10679;
assign n_10681 = ~x_263 & ~n_10680;
assign n_10682 =  x_263 & ~n_10679;
assign n_10683 = ~n_10678 &  n_10682;
assign n_10684 =  n_10522 & ~n_10683;
assign n_10685 = ~n_10681 &  n_10684;
assign n_10686 = ~n_10673 & ~n_10685;
assign n_10687 =  n_10661 &  n_10686;
assign n_10688 =  x_1095 & ~n_10687;
assign n_10689 = ~x_1095 &  n_10687;
assign n_10690 = ~n_10688 & ~n_10689;
assign n_10691 = ~x_1702 &  n_10674;
assign n_10692 =  x_1702 & ~n_10674;
assign n_10693 = ~n_10691 & ~n_10692;
assign n_10694 = ~n_10678 & ~n_10682;
assign n_10695 =  n_10693 & ~n_10694;
assign n_10696 = ~n_10693 &  n_10694;
assign n_10697 = ~n_10695 & ~n_10696;
assign n_10698 = ~x_262 & ~n_10697;
assign n_10699 =  x_262 & ~n_10696;
assign n_10700 = ~n_10695 &  n_10699;
assign n_10701 =  n_10522 & ~n_10700;
assign n_10702 = ~n_10698 &  n_10701;
assign n_10703 =  x_1094 &  n_10525;
assign n_10704 = ~x_870 &  n_10656;
assign n_10705 =  x_870 & ~n_10656;
assign n_10706 = ~n_10704 & ~n_10705;
assign n_10707 =  n_10517 &  n_10706;
assign n_10708 = ~n_10703 & ~n_10707;
assign n_10709 = ~n_10702 &  n_10708;
assign n_10710 = ~x_2342 &  n_10662;
assign n_10711 =  x_2342 & ~n_10662;
assign n_10712 = ~n_10710 & ~n_10711;
assign n_10713 = ~n_10666 & ~n_10670;
assign n_10714 =  n_10712 & ~n_10713;
assign n_10715 = ~n_10712 &  n_10713;
assign n_10716 = ~n_10714 & ~n_10715;
assign n_10717 = ~x_454 & ~n_10716;
assign n_10718 =  x_454 & ~n_10715;
assign n_10719 = ~n_10714 &  n_10718;
assign n_10720 =  n_10523 & ~n_10719;
assign n_10721 = ~n_10717 &  n_10720;
assign n_10722 = ~x_230 &  n_10643;
assign n_10723 =  x_230 & ~n_10643;
assign n_10724 = ~n_10722 & ~n_10723;
assign n_10725 = ~n_10647 & ~n_10651;
assign n_10726 =  n_10724 & ~n_10725;
assign n_10727 = ~n_10724 &  n_10725;
assign n_10728 = ~n_10726 & ~n_10727;
assign n_10729 = ~x_2694 & ~n_10728;
assign n_10730 =  x_2694 & ~n_10727;
assign n_10731 = ~n_10726 &  n_10730;
assign n_10732 =  n_10519 & ~n_10731;
assign n_10733 = ~n_10729 &  n_10732;
assign n_10734 = ~n_10721 & ~n_10733;
assign n_10735 =  n_10709 &  n_10734;
assign n_10736 =  x_1094 & ~n_10735;
assign n_10737 = ~x_1094 &  n_10735;
assign n_10738 = ~n_10736 & ~n_10737;
assign n_10739 = ~x_1701 &  n_10691;
assign n_10740 =  x_1701 & ~n_10691;
assign n_10741 = ~n_10739 & ~n_10740;
assign n_10742 = ~n_10695 & ~n_10699;
assign n_10743 =  n_10741 & ~n_10742;
assign n_10744 = ~n_10741 &  n_10742;
assign n_10745 = ~n_10743 & ~n_10744;
assign n_10746 = ~x_261 & ~n_10745;
assign n_10747 =  x_261 & ~n_10744;
assign n_10748 = ~n_10743 &  n_10747;
assign n_10749 =  n_10522 & ~n_10748;
assign n_10750 = ~n_10746 &  n_10749;
assign n_10751 =  x_1093 &  n_10525;
assign n_10752 = ~x_869 &  n_10704;
assign n_10753 =  x_869 & ~n_10704;
assign n_10754 = ~n_10752 & ~n_10753;
assign n_10755 =  n_10517 &  n_10754;
assign n_10756 = ~n_10751 & ~n_10755;
assign n_10757 = ~n_10750 &  n_10756;
assign n_10758 = ~x_2341 &  n_10710;
assign n_10759 =  x_2341 & ~n_10710;
assign n_10760 = ~n_10758 & ~n_10759;
assign n_10761 = ~n_10714 & ~n_10718;
assign n_10762 =  n_10760 & ~n_10761;
assign n_10763 = ~n_10760 &  n_10761;
assign n_10764 = ~n_10762 & ~n_10763;
assign n_10765 = ~x_453 & ~n_10764;
assign n_10766 =  x_453 & ~n_10763;
assign n_10767 = ~n_10762 &  n_10766;
assign n_10768 =  n_10523 & ~n_10767;
assign n_10769 = ~n_10765 &  n_10768;
assign n_10770 = ~x_229 &  n_10722;
assign n_10771 =  x_229 & ~n_10722;
assign n_10772 = ~n_10770 & ~n_10771;
assign n_10773 = ~n_10726 & ~n_10730;
assign n_10774 =  n_10772 & ~n_10773;
assign n_10775 = ~n_10772 &  n_10773;
assign n_10776 = ~n_10774 & ~n_10775;
assign n_10777 = ~x_2693 & ~n_10776;
assign n_10778 =  x_2693 & ~n_10775;
assign n_10779 = ~n_10774 &  n_10778;
assign n_10780 =  n_10519 & ~n_10779;
assign n_10781 = ~n_10777 &  n_10780;
assign n_10782 = ~n_10769 & ~n_10781;
assign n_10783 =  n_10757 &  n_10782;
assign n_10784 =  x_1093 & ~n_10783;
assign n_10785 = ~x_1093 &  n_10783;
assign n_10786 = ~n_10784 & ~n_10785;
assign n_10787 = ~x_1700 &  n_10739;
assign n_10788 =  x_1700 & ~n_10739;
assign n_10789 = ~n_10787 & ~n_10788;
assign n_10790 = ~n_10743 & ~n_10747;
assign n_10791 =  n_10789 & ~n_10790;
assign n_10792 = ~n_10789 &  n_10790;
assign n_10793 = ~n_10791 & ~n_10792;
assign n_10794 = ~x_260 & ~n_10793;
assign n_10795 =  x_260 & ~n_10792;
assign n_10796 = ~n_10791 &  n_10795;
assign n_10797 =  n_10522 & ~n_10796;
assign n_10798 = ~n_10794 &  n_10797;
assign n_10799 =  x_1092 &  n_10525;
assign n_10800 =  x_868 & ~n_10752;
assign n_10801 = ~x_868 &  n_10752;
assign n_10802 =  n_10517 & ~n_10801;
assign n_10803 = ~n_10800 &  n_10802;
assign n_10804 = ~n_10799 & ~n_10803;
assign n_10805 = ~n_10798 &  n_10804;
assign n_10806 = ~x_2340 &  n_10758;
assign n_10807 =  x_2340 & ~n_10758;
assign n_10808 = ~n_10806 & ~n_10807;
assign n_10809 = ~n_10762 & ~n_10766;
assign n_10810 =  n_10808 & ~n_10809;
assign n_10811 = ~n_10808 &  n_10809;
assign n_10812 = ~n_10810 & ~n_10811;
assign n_10813 = ~x_452 & ~n_10812;
assign n_10814 =  x_452 & ~n_10811;
assign n_10815 = ~n_10810 &  n_10814;
assign n_10816 =  n_10523 & ~n_10815;
assign n_10817 = ~n_10813 &  n_10816;
assign n_10818 = ~x_228 &  n_10770;
assign n_10819 =  x_228 & ~n_10770;
assign n_10820 = ~n_10818 & ~n_10819;
assign n_10821 = ~n_10774 & ~n_10778;
assign n_10822 =  n_10820 & ~n_10821;
assign n_10823 = ~n_10820 &  n_10821;
assign n_10824 = ~n_10822 & ~n_10823;
assign n_10825 = ~x_2692 & ~n_10824;
assign n_10826 =  x_2692 & ~n_10823;
assign n_10827 = ~n_10822 &  n_10826;
assign n_10828 =  n_10519 & ~n_10827;
assign n_10829 = ~n_10825 &  n_10828;
assign n_10830 = ~n_10817 & ~n_10829;
assign n_10831 =  n_10805 &  n_10830;
assign n_10832 =  x_1092 & ~n_10831;
assign n_10833 = ~x_1092 &  n_10831;
assign n_10834 = ~n_10832 & ~n_10833;
assign n_10835 = ~x_1699 &  n_10787;
assign n_10836 =  x_1699 & ~n_10787;
assign n_10837 = ~n_10835 & ~n_10836;
assign n_10838 = ~n_10791 & ~n_10795;
assign n_10839 =  n_10837 & ~n_10838;
assign n_10840 = ~n_10837 &  n_10838;
assign n_10841 = ~n_10839 & ~n_10840;
assign n_10842 = ~x_259 & ~n_10841;
assign n_10843 =  x_259 & ~n_10840;
assign n_10844 = ~n_10839 &  n_10843;
assign n_10845 =  n_10522 & ~n_10844;
assign n_10846 = ~n_10842 &  n_10845;
assign n_10847 =  x_1091 &  n_10525;
assign n_10848 =  x_867 & ~n_10801;
assign n_10849 = ~x_867 &  n_10801;
assign n_10850 =  n_10517 & ~n_10849;
assign n_10851 = ~n_10848 &  n_10850;
assign n_10852 = ~n_10847 & ~n_10851;
assign n_10853 = ~n_10846 &  n_10852;
assign n_10854 = ~x_2339 &  n_10806;
assign n_10855 =  x_2339 & ~n_10806;
assign n_10856 = ~n_10854 & ~n_10855;
assign n_10857 = ~n_10810 & ~n_10814;
assign n_10858 =  n_10856 & ~n_10857;
assign n_10859 = ~n_10856 &  n_10857;
assign n_10860 = ~n_10858 & ~n_10859;
assign n_10861 = ~x_451 & ~n_10860;
assign n_10862 =  x_451 & ~n_10859;
assign n_10863 = ~n_10858 &  n_10862;
assign n_10864 =  n_10523 & ~n_10863;
assign n_10865 = ~n_10861 &  n_10864;
assign n_10866 = ~x_227 &  n_10818;
assign n_10867 =  x_227 & ~n_10818;
assign n_10868 = ~n_10866 & ~n_10867;
assign n_10869 = ~n_10822 & ~n_10826;
assign n_10870 =  n_10868 & ~n_10869;
assign n_10871 = ~n_10868 &  n_10869;
assign n_10872 = ~n_10870 & ~n_10871;
assign n_10873 = ~x_2691 & ~n_10872;
assign n_10874 =  x_2691 & ~n_10871;
assign n_10875 = ~n_10870 &  n_10874;
assign n_10876 =  n_10519 & ~n_10875;
assign n_10877 = ~n_10873 &  n_10876;
assign n_10878 = ~n_10865 & ~n_10877;
assign n_10879 =  n_10853 &  n_10878;
assign n_10880 =  x_1091 & ~n_10879;
assign n_10881 = ~x_1091 &  n_10879;
assign n_10882 = ~n_10880 & ~n_10881;
assign n_10883 = ~x_1698 &  n_10835;
assign n_10884 =  x_1698 & ~n_10835;
assign n_10885 = ~n_10883 & ~n_10884;
assign n_10886 = ~n_10839 & ~n_10843;
assign n_10887 =  n_10885 & ~n_10886;
assign n_10888 = ~n_10885 &  n_10886;
assign n_10889 = ~n_10887 & ~n_10888;
assign n_10890 = ~x_258 & ~n_10889;
assign n_10891 =  x_258 & ~n_10888;
assign n_10892 = ~n_10887 &  n_10891;
assign n_10893 =  n_10522 & ~n_10892;
assign n_10894 = ~n_10890 &  n_10893;
assign n_10895 =  x_1090 &  n_10525;
assign n_10896 =  x_866 & ~n_10849;
assign n_10897 = ~x_866 &  n_10849;
assign n_10898 =  n_10517 & ~n_10897;
assign n_10899 = ~n_10896 &  n_10898;
assign n_10900 = ~n_10895 & ~n_10899;
assign n_10901 = ~n_10894 &  n_10900;
assign n_10902 = ~x_2338 &  n_10854;
assign n_10903 =  x_2338 & ~n_10854;
assign n_10904 = ~n_10902 & ~n_10903;
assign n_10905 = ~n_10858 & ~n_10862;
assign n_10906 =  n_10904 & ~n_10905;
assign n_10907 = ~n_10904 &  n_10905;
assign n_10908 = ~n_10906 & ~n_10907;
assign n_10909 = ~x_450 & ~n_10908;
assign n_10910 =  x_450 & ~n_10907;
assign n_10911 = ~n_10906 &  n_10910;
assign n_10912 =  n_10523 & ~n_10911;
assign n_10913 = ~n_10909 &  n_10912;
assign n_10914 = ~x_226 &  n_10866;
assign n_10915 =  x_226 & ~n_10866;
assign n_10916 = ~n_10914 & ~n_10915;
assign n_10917 = ~n_10870 & ~n_10874;
assign n_10918 =  n_10916 & ~n_10917;
assign n_10919 = ~n_10916 &  n_10917;
assign n_10920 = ~n_10918 & ~n_10919;
assign n_10921 = ~x_2690 & ~n_10920;
assign n_10922 =  x_2690 & ~n_10919;
assign n_10923 = ~n_10918 &  n_10922;
assign n_10924 =  n_10519 & ~n_10923;
assign n_10925 = ~n_10921 &  n_10924;
assign n_10926 = ~n_10913 & ~n_10925;
assign n_10927 =  n_10901 &  n_10926;
assign n_10928 =  x_1090 & ~n_10927;
assign n_10929 = ~x_1090 &  n_10927;
assign n_10930 = ~n_10928 & ~n_10929;
assign n_10931 = ~x_1697 &  n_10883;
assign n_10932 =  x_1697 & ~n_10883;
assign n_10933 = ~n_10931 & ~n_10932;
assign n_10934 = ~n_10887 & ~n_10891;
assign n_10935 =  n_10933 & ~n_10934;
assign n_10936 = ~n_10933 &  n_10934;
assign n_10937 = ~n_10935 & ~n_10936;
assign n_10938 = ~x_257 & ~n_10937;
assign n_10939 =  x_257 & ~n_10936;
assign n_10940 = ~n_10935 &  n_10939;
assign n_10941 =  n_10522 & ~n_10940;
assign n_10942 = ~n_10938 &  n_10941;
assign n_10943 =  x_1089 &  n_10525;
assign n_10944 =  x_865 & ~n_10897;
assign n_10945 = ~x_865 &  n_10897;
assign n_10946 =  n_10517 & ~n_10945;
assign n_10947 = ~n_10944 &  n_10946;
assign n_10948 = ~n_10943 & ~n_10947;
assign n_10949 = ~n_10942 &  n_10948;
assign n_10950 = ~x_2337 &  n_10902;
assign n_10951 =  x_2337 & ~n_10902;
assign n_10952 = ~n_10950 & ~n_10951;
assign n_10953 = ~n_10906 & ~n_10910;
assign n_10954 =  n_10952 & ~n_10953;
assign n_10955 = ~n_10952 &  n_10953;
assign n_10956 = ~n_10954 & ~n_10955;
assign n_10957 = ~x_449 & ~n_10956;
assign n_10958 =  x_449 & ~n_10955;
assign n_10959 = ~n_10954 &  n_10958;
assign n_10960 =  n_10523 & ~n_10959;
assign n_10961 = ~n_10957 &  n_10960;
assign n_10962 = ~x_225 &  n_10914;
assign n_10963 =  x_225 & ~n_10914;
assign n_10964 = ~n_10962 & ~n_10963;
assign n_10965 = ~n_10918 & ~n_10922;
assign n_10966 =  n_10964 & ~n_10965;
assign n_10967 = ~n_10964 &  n_10965;
assign n_10968 = ~n_10966 & ~n_10967;
assign n_10969 = ~x_2689 & ~n_10968;
assign n_10970 =  x_2689 & ~n_10967;
assign n_10971 = ~n_10966 &  n_10970;
assign n_10972 =  n_10519 & ~n_10971;
assign n_10973 = ~n_10969 &  n_10972;
assign n_10974 = ~n_10961 & ~n_10973;
assign n_10975 =  n_10949 &  n_10974;
assign n_10976 =  x_1089 & ~n_10975;
assign n_10977 = ~x_1089 &  n_10975;
assign n_10978 = ~n_10976 & ~n_10977;
assign n_10979 = ~x_1696 &  n_10931;
assign n_10980 =  x_1696 & ~n_10931;
assign n_10981 = ~n_10979 & ~n_10980;
assign n_10982 = ~n_10935 & ~n_10939;
assign n_10983 =  n_10981 & ~n_10982;
assign n_10984 = ~n_10981 &  n_10982;
assign n_10985 = ~n_10983 & ~n_10984;
assign n_10986 = ~x_256 & ~n_10985;
assign n_10987 =  x_256 & ~n_10984;
assign n_10988 = ~n_10983 &  n_10987;
assign n_10989 =  n_10522 & ~n_10988;
assign n_10990 = ~n_10986 &  n_10989;
assign n_10991 =  x_1088 &  n_10525;
assign n_10992 =  x_864 & ~n_10945;
assign n_10993 = ~x_864 &  n_10945;
assign n_10994 =  n_10517 & ~n_10993;
assign n_10995 = ~n_10992 &  n_10994;
assign n_10996 = ~n_10991 & ~n_10995;
assign n_10997 = ~n_10990 &  n_10996;
assign n_10998 = ~x_2336 &  n_10950;
assign n_10999 =  x_2336 & ~n_10950;
assign n_11000 = ~n_10998 & ~n_10999;
assign n_11001 = ~n_10954 & ~n_10958;
assign n_11002 =  n_11000 & ~n_11001;
assign n_11003 = ~n_11000 &  n_11001;
assign n_11004 = ~n_11002 & ~n_11003;
assign n_11005 = ~x_448 & ~n_11004;
assign n_11006 =  x_448 & ~n_11003;
assign n_11007 = ~n_11002 &  n_11006;
assign n_11008 =  n_10523 & ~n_11007;
assign n_11009 = ~n_11005 &  n_11008;
assign n_11010 = ~x_224 &  n_10962;
assign n_11011 =  x_224 & ~n_10962;
assign n_11012 = ~n_11010 & ~n_11011;
assign n_11013 = ~n_10966 & ~n_10970;
assign n_11014 =  n_11012 & ~n_11013;
assign n_11015 = ~n_11012 &  n_11013;
assign n_11016 = ~n_11014 & ~n_11015;
assign n_11017 = ~x_2688 & ~n_11016;
assign n_11018 =  x_2688 & ~n_11015;
assign n_11019 = ~n_11014 &  n_11018;
assign n_11020 =  n_10519 & ~n_11019;
assign n_11021 = ~n_11017 &  n_11020;
assign n_11022 = ~n_11009 & ~n_11021;
assign n_11023 =  n_10997 &  n_11022;
assign n_11024 =  x_1088 & ~n_11023;
assign n_11025 = ~x_1088 &  n_11023;
assign n_11026 = ~n_11024 & ~n_11025;
assign n_11027 = ~x_1695 &  n_10979;
assign n_11028 =  x_1695 & ~n_10979;
assign n_11029 = ~n_11027 & ~n_11028;
assign n_11030 = ~n_10983 & ~n_10987;
assign n_11031 =  n_11029 & ~n_11030;
assign n_11032 = ~n_11029 &  n_11030;
assign n_11033 = ~n_11031 & ~n_11032;
assign n_11034 = ~x_255 & ~n_11033;
assign n_11035 =  x_255 & ~n_11032;
assign n_11036 = ~n_11031 &  n_11035;
assign n_11037 =  n_10522 & ~n_11036;
assign n_11038 = ~n_11034 &  n_11037;
assign n_11039 =  x_1087 &  n_10525;
assign n_11040 =  x_863 & ~n_10993;
assign n_11041 = ~x_863 &  n_10993;
assign n_11042 =  n_10517 & ~n_11041;
assign n_11043 = ~n_11040 &  n_11042;
assign n_11044 = ~n_11039 & ~n_11043;
assign n_11045 = ~n_11038 &  n_11044;
assign n_11046 = ~x_2335 &  n_10998;
assign n_11047 =  x_2335 & ~n_10998;
assign n_11048 = ~n_11046 & ~n_11047;
assign n_11049 = ~n_11002 & ~n_11006;
assign n_11050 =  n_11048 & ~n_11049;
assign n_11051 = ~n_11048 &  n_11049;
assign n_11052 = ~n_11050 & ~n_11051;
assign n_11053 = ~x_447 & ~n_11052;
assign n_11054 =  x_447 & ~n_11051;
assign n_11055 = ~n_11050 &  n_11054;
assign n_11056 =  n_10523 & ~n_11055;
assign n_11057 = ~n_11053 &  n_11056;
assign n_11058 = ~x_223 &  n_11010;
assign n_11059 =  x_223 & ~n_11010;
assign n_11060 = ~n_11058 & ~n_11059;
assign n_11061 = ~n_11014 & ~n_11018;
assign n_11062 =  n_11060 & ~n_11061;
assign n_11063 = ~n_11060 &  n_11061;
assign n_11064 = ~n_11062 & ~n_11063;
assign n_11065 = ~x_2687 & ~n_11064;
assign n_11066 =  x_2687 & ~n_11063;
assign n_11067 = ~n_11062 &  n_11066;
assign n_11068 =  n_10519 & ~n_11067;
assign n_11069 = ~n_11065 &  n_11068;
assign n_11070 = ~n_11057 & ~n_11069;
assign n_11071 =  n_11045 &  n_11070;
assign n_11072 =  x_1087 & ~n_11071;
assign n_11073 = ~x_1087 &  n_11071;
assign n_11074 = ~n_11072 & ~n_11073;
assign n_11075 = ~x_1694 &  n_11027;
assign n_11076 =  x_1694 & ~n_11027;
assign n_11077 = ~n_11075 & ~n_11076;
assign n_11078 = ~n_11031 & ~n_11035;
assign n_11079 =  n_11077 & ~n_11078;
assign n_11080 = ~n_11077 &  n_11078;
assign n_11081 = ~n_11079 & ~n_11080;
assign n_11082 = ~x_254 & ~n_11081;
assign n_11083 =  x_254 & ~n_11080;
assign n_11084 = ~n_11079 &  n_11083;
assign n_11085 =  n_10522 & ~n_11084;
assign n_11086 = ~n_11082 &  n_11085;
assign n_11087 =  x_1086 &  n_10525;
assign n_11088 =  x_862 & ~n_11041;
assign n_11089 = ~x_862 &  n_11041;
assign n_11090 =  n_10517 & ~n_11089;
assign n_11091 = ~n_11088 &  n_11090;
assign n_11092 = ~n_11087 & ~n_11091;
assign n_11093 = ~n_11086 &  n_11092;
assign n_11094 = ~x_2334 &  n_11046;
assign n_11095 =  x_2334 & ~n_11046;
assign n_11096 = ~n_11094 & ~n_11095;
assign n_11097 = ~n_11050 & ~n_11054;
assign n_11098 =  n_11096 & ~n_11097;
assign n_11099 = ~n_11096 &  n_11097;
assign n_11100 = ~n_11098 & ~n_11099;
assign n_11101 = ~x_446 & ~n_11100;
assign n_11102 =  x_446 & ~n_11099;
assign n_11103 = ~n_11098 &  n_11102;
assign n_11104 =  n_10523 & ~n_11103;
assign n_11105 = ~n_11101 &  n_11104;
assign n_11106 = ~x_222 &  n_11058;
assign n_11107 =  x_222 & ~n_11058;
assign n_11108 = ~n_11106 & ~n_11107;
assign n_11109 = ~n_11062 & ~n_11066;
assign n_11110 =  n_11108 & ~n_11109;
assign n_11111 = ~n_11108 &  n_11109;
assign n_11112 = ~n_11110 & ~n_11111;
assign n_11113 = ~x_2686 & ~n_11112;
assign n_11114 =  x_2686 & ~n_11111;
assign n_11115 = ~n_11110 &  n_11114;
assign n_11116 =  n_10519 & ~n_11115;
assign n_11117 = ~n_11113 &  n_11116;
assign n_11118 = ~n_11105 & ~n_11117;
assign n_11119 =  n_11093 &  n_11118;
assign n_11120 =  x_1086 & ~n_11119;
assign n_11121 = ~x_1086 &  n_11119;
assign n_11122 = ~n_11120 & ~n_11121;
assign n_11123 = ~x_1693 &  n_11075;
assign n_11124 =  x_1693 & ~n_11075;
assign n_11125 = ~n_11123 & ~n_11124;
assign n_11126 = ~n_11079 & ~n_11083;
assign n_11127 =  n_11125 & ~n_11126;
assign n_11128 = ~n_11125 &  n_11126;
assign n_11129 = ~n_11127 & ~n_11128;
assign n_11130 = ~x_253 & ~n_11129;
assign n_11131 =  x_253 & ~n_11128;
assign n_11132 = ~n_11127 &  n_11131;
assign n_11133 =  n_10522 & ~n_11132;
assign n_11134 = ~n_11130 &  n_11133;
assign n_11135 =  x_1085 &  n_10525;
assign n_11136 =  x_861 & ~n_11089;
assign n_11137 = ~x_861 &  n_11089;
assign n_11138 =  n_10517 & ~n_11137;
assign n_11139 = ~n_11136 &  n_11138;
assign n_11140 = ~n_11135 & ~n_11139;
assign n_11141 = ~n_11134 &  n_11140;
assign n_11142 = ~x_2333 &  n_11094;
assign n_11143 =  x_2333 & ~n_11094;
assign n_11144 = ~n_11142 & ~n_11143;
assign n_11145 = ~n_11098 & ~n_11102;
assign n_11146 =  n_11144 & ~n_11145;
assign n_11147 = ~n_11144 &  n_11145;
assign n_11148 = ~n_11146 & ~n_11147;
assign n_11149 = ~x_445 & ~n_11148;
assign n_11150 =  x_445 & ~n_11147;
assign n_11151 = ~n_11146 &  n_11150;
assign n_11152 =  n_10523 & ~n_11151;
assign n_11153 = ~n_11149 &  n_11152;
assign n_11154 = ~x_221 &  n_11106;
assign n_11155 =  x_221 & ~n_11106;
assign n_11156 = ~n_11154 & ~n_11155;
assign n_11157 = ~n_11110 & ~n_11114;
assign n_11158 =  n_11156 & ~n_11157;
assign n_11159 = ~n_11156 &  n_11157;
assign n_11160 = ~n_11158 & ~n_11159;
assign n_11161 = ~x_2685 & ~n_11160;
assign n_11162 =  x_2685 & ~n_11159;
assign n_11163 = ~n_11158 &  n_11162;
assign n_11164 =  n_10519 & ~n_11163;
assign n_11165 = ~n_11161 &  n_11164;
assign n_11166 = ~n_11153 & ~n_11165;
assign n_11167 =  n_11141 &  n_11166;
assign n_11168 =  x_1085 & ~n_11167;
assign n_11169 = ~x_1085 &  n_11167;
assign n_11170 = ~n_11168 & ~n_11169;
assign n_11171 = ~x_1692 &  n_11123;
assign n_11172 =  x_1692 & ~n_11123;
assign n_11173 = ~n_11171 & ~n_11172;
assign n_11174 = ~n_11127 & ~n_11131;
assign n_11175 =  n_11173 & ~n_11174;
assign n_11176 = ~n_11173 &  n_11174;
assign n_11177 = ~n_11175 & ~n_11176;
assign n_11178 = ~x_252 & ~n_11177;
assign n_11179 =  x_252 & ~n_11176;
assign n_11180 = ~n_11175 &  n_11179;
assign n_11181 =  n_10522 & ~n_11180;
assign n_11182 = ~n_11178 &  n_11181;
assign n_11183 =  x_1084 &  n_10525;
assign n_11184 =  x_860 & ~n_11137;
assign n_11185 = ~x_860 &  n_11137;
assign n_11186 =  n_10517 & ~n_11185;
assign n_11187 = ~n_11184 &  n_11186;
assign n_11188 = ~n_11183 & ~n_11187;
assign n_11189 = ~n_11182 &  n_11188;
assign n_11190 = ~x_2332 &  n_11142;
assign n_11191 =  x_2332 & ~n_11142;
assign n_11192 = ~n_11190 & ~n_11191;
assign n_11193 = ~n_11146 & ~n_11150;
assign n_11194 =  n_11192 & ~n_11193;
assign n_11195 = ~n_11192 &  n_11193;
assign n_11196 = ~n_11194 & ~n_11195;
assign n_11197 = ~x_444 & ~n_11196;
assign n_11198 =  x_444 & ~n_11195;
assign n_11199 = ~n_11194 &  n_11198;
assign n_11200 =  n_10523 & ~n_11199;
assign n_11201 = ~n_11197 &  n_11200;
assign n_11202 = ~x_220 &  n_11154;
assign n_11203 =  x_220 & ~n_11154;
assign n_11204 = ~n_11202 & ~n_11203;
assign n_11205 = ~n_11158 & ~n_11162;
assign n_11206 =  n_11204 & ~n_11205;
assign n_11207 = ~n_11204 &  n_11205;
assign n_11208 = ~n_11206 & ~n_11207;
assign n_11209 = ~x_2684 & ~n_11208;
assign n_11210 =  x_2684 & ~n_11207;
assign n_11211 = ~n_11206 &  n_11210;
assign n_11212 =  n_10519 & ~n_11211;
assign n_11213 = ~n_11209 &  n_11212;
assign n_11214 = ~n_11201 & ~n_11213;
assign n_11215 =  n_11189 &  n_11214;
assign n_11216 =  x_1084 & ~n_11215;
assign n_11217 = ~x_1084 &  n_11215;
assign n_11218 = ~n_11216 & ~n_11217;
assign n_11219 = ~x_1691 &  n_11171;
assign n_11220 =  x_1691 & ~n_11171;
assign n_11221 = ~n_11219 & ~n_11220;
assign n_11222 = ~n_11175 & ~n_11179;
assign n_11223 =  n_11221 & ~n_11222;
assign n_11224 = ~n_11221 &  n_11222;
assign n_11225 = ~n_11223 & ~n_11224;
assign n_11226 = ~x_251 & ~n_11225;
assign n_11227 =  x_251 & ~n_11224;
assign n_11228 = ~n_11223 &  n_11227;
assign n_11229 =  n_10522 & ~n_11228;
assign n_11230 = ~n_11226 &  n_11229;
assign n_11231 =  x_1083 &  n_10525;
assign n_11232 =  x_859 & ~n_11185;
assign n_11233 = ~x_859 &  n_11185;
assign n_11234 =  n_10517 & ~n_11233;
assign n_11235 = ~n_11232 &  n_11234;
assign n_11236 = ~n_11231 & ~n_11235;
assign n_11237 = ~n_11230 &  n_11236;
assign n_11238 = ~x_2331 &  n_11190;
assign n_11239 =  x_2331 & ~n_11190;
assign n_11240 = ~n_11238 & ~n_11239;
assign n_11241 = ~n_11194 & ~n_11198;
assign n_11242 =  n_11240 & ~n_11241;
assign n_11243 = ~n_11240 &  n_11241;
assign n_11244 = ~n_11242 & ~n_11243;
assign n_11245 = ~x_443 & ~n_11244;
assign n_11246 =  x_443 & ~n_11243;
assign n_11247 = ~n_11242 &  n_11246;
assign n_11248 =  n_10523 & ~n_11247;
assign n_11249 = ~n_11245 &  n_11248;
assign n_11250 = ~x_219 &  n_11202;
assign n_11251 =  x_219 & ~n_11202;
assign n_11252 = ~n_11250 & ~n_11251;
assign n_11253 = ~n_11206 & ~n_11210;
assign n_11254 =  n_11252 & ~n_11253;
assign n_11255 = ~n_11252 &  n_11253;
assign n_11256 = ~n_11254 & ~n_11255;
assign n_11257 = ~x_2683 & ~n_11256;
assign n_11258 =  x_2683 & ~n_11255;
assign n_11259 = ~n_11254 &  n_11258;
assign n_11260 =  n_10519 & ~n_11259;
assign n_11261 = ~n_11257 &  n_11260;
assign n_11262 = ~n_11249 & ~n_11261;
assign n_11263 =  n_11237 &  n_11262;
assign n_11264 =  x_1083 & ~n_11263;
assign n_11265 = ~x_1083 &  n_11263;
assign n_11266 = ~n_11264 & ~n_11265;
assign n_11267 = ~x_1690 &  n_11219;
assign n_11268 =  x_1690 & ~n_11219;
assign n_11269 = ~n_11267 & ~n_11268;
assign n_11270 = ~n_11223 & ~n_11227;
assign n_11271 =  n_11269 & ~n_11270;
assign n_11272 = ~n_11269 &  n_11270;
assign n_11273 = ~n_11271 & ~n_11272;
assign n_11274 = ~x_250 & ~n_11273;
assign n_11275 =  x_250 & ~n_11272;
assign n_11276 = ~n_11271 &  n_11275;
assign n_11277 =  n_10522 & ~n_11276;
assign n_11278 = ~n_11274 &  n_11277;
assign n_11279 =  x_1082 &  n_10525;
assign n_11280 =  x_858 & ~n_11233;
assign n_11281 = ~x_858 &  n_11233;
assign n_11282 =  n_10517 & ~n_11281;
assign n_11283 = ~n_11280 &  n_11282;
assign n_11284 = ~n_11279 & ~n_11283;
assign n_11285 = ~n_11278 &  n_11284;
assign n_11286 = ~x_2330 &  n_11238;
assign n_11287 =  x_2330 & ~n_11238;
assign n_11288 = ~n_11286 & ~n_11287;
assign n_11289 = ~n_11242 & ~n_11246;
assign n_11290 =  n_11288 & ~n_11289;
assign n_11291 = ~n_11288 &  n_11289;
assign n_11292 = ~n_11290 & ~n_11291;
assign n_11293 = ~x_442 & ~n_11292;
assign n_11294 =  x_442 & ~n_11291;
assign n_11295 = ~n_11290 &  n_11294;
assign n_11296 =  n_10523 & ~n_11295;
assign n_11297 = ~n_11293 &  n_11296;
assign n_11298 = ~x_218 &  n_11250;
assign n_11299 =  x_218 & ~n_11250;
assign n_11300 = ~n_11298 & ~n_11299;
assign n_11301 = ~n_11254 & ~n_11258;
assign n_11302 =  n_11300 & ~n_11301;
assign n_11303 = ~n_11300 &  n_11301;
assign n_11304 = ~n_11302 & ~n_11303;
assign n_11305 = ~x_2682 & ~n_11304;
assign n_11306 =  x_2682 & ~n_11303;
assign n_11307 = ~n_11302 &  n_11306;
assign n_11308 =  n_10519 & ~n_11307;
assign n_11309 = ~n_11305 &  n_11308;
assign n_11310 = ~n_11297 & ~n_11309;
assign n_11311 =  n_11285 &  n_11310;
assign n_11312 =  x_1082 & ~n_11311;
assign n_11313 = ~x_1082 &  n_11311;
assign n_11314 = ~n_11312 & ~n_11313;
assign n_11315 = ~x_1689 &  n_11267;
assign n_11316 =  x_1689 & ~n_11267;
assign n_11317 = ~n_11315 & ~n_11316;
assign n_11318 = ~n_11271 & ~n_11275;
assign n_11319 =  n_11317 & ~n_11318;
assign n_11320 = ~n_11317 &  n_11318;
assign n_11321 = ~n_11319 & ~n_11320;
assign n_11322 = ~x_249 & ~n_11321;
assign n_11323 =  x_249 & ~n_11320;
assign n_11324 = ~n_11319 &  n_11323;
assign n_11325 =  n_10522 & ~n_11324;
assign n_11326 = ~n_11322 &  n_11325;
assign n_11327 =  x_1081 &  n_10525;
assign n_11328 =  x_857 & ~n_11281;
assign n_11329 = ~x_857 &  n_11281;
assign n_11330 =  n_10517 & ~n_11329;
assign n_11331 = ~n_11328 &  n_11330;
assign n_11332 = ~n_11327 & ~n_11331;
assign n_11333 = ~n_11326 &  n_11332;
assign n_11334 = ~x_2329 &  n_11286;
assign n_11335 =  x_2329 & ~n_11286;
assign n_11336 = ~n_11334 & ~n_11335;
assign n_11337 = ~n_11290 & ~n_11294;
assign n_11338 =  n_11336 & ~n_11337;
assign n_11339 = ~n_11336 &  n_11337;
assign n_11340 = ~n_11338 & ~n_11339;
assign n_11341 = ~x_441 & ~n_11340;
assign n_11342 =  x_441 & ~n_11339;
assign n_11343 = ~n_11338 &  n_11342;
assign n_11344 =  n_10523 & ~n_11343;
assign n_11345 = ~n_11341 &  n_11344;
assign n_11346 = ~x_217 &  n_11298;
assign n_11347 =  x_217 & ~n_11298;
assign n_11348 = ~n_11346 & ~n_11347;
assign n_11349 = ~n_11302 & ~n_11306;
assign n_11350 =  n_11348 & ~n_11349;
assign n_11351 = ~n_11348 &  n_11349;
assign n_11352 = ~n_11350 & ~n_11351;
assign n_11353 = ~x_2681 & ~n_11352;
assign n_11354 =  x_2681 & ~n_11351;
assign n_11355 = ~n_11350 &  n_11354;
assign n_11356 =  n_10519 & ~n_11355;
assign n_11357 = ~n_11353 &  n_11356;
assign n_11358 = ~n_11345 & ~n_11357;
assign n_11359 =  n_11333 &  n_11358;
assign n_11360 =  x_1081 & ~n_11359;
assign n_11361 = ~x_1081 &  n_11359;
assign n_11362 = ~n_11360 & ~n_11361;
assign n_11363 = ~x_1688 &  n_11315;
assign n_11364 =  x_1688 & ~n_11315;
assign n_11365 = ~n_11363 & ~n_11364;
assign n_11366 = ~n_11319 & ~n_11323;
assign n_11367 =  n_11365 & ~n_11366;
assign n_11368 = ~n_11365 &  n_11366;
assign n_11369 = ~n_11367 & ~n_11368;
assign n_11370 = ~x_248 & ~n_11369;
assign n_11371 =  x_248 & ~n_11368;
assign n_11372 = ~n_11367 &  n_11371;
assign n_11373 =  n_10522 & ~n_11372;
assign n_11374 = ~n_11370 &  n_11373;
assign n_11375 =  x_1080 &  n_10525;
assign n_11376 =  x_856 & ~n_11329;
assign n_11377 = ~x_856 &  n_11329;
assign n_11378 =  n_10517 & ~n_11377;
assign n_11379 = ~n_11376 &  n_11378;
assign n_11380 = ~n_11375 & ~n_11379;
assign n_11381 = ~n_11374 &  n_11380;
assign n_11382 = ~x_2328 &  n_11334;
assign n_11383 =  x_2328 & ~n_11334;
assign n_11384 = ~n_11382 & ~n_11383;
assign n_11385 = ~n_11338 & ~n_11342;
assign n_11386 =  n_11384 & ~n_11385;
assign n_11387 = ~n_11384 &  n_11385;
assign n_11388 = ~n_11386 & ~n_11387;
assign n_11389 = ~x_440 & ~n_11388;
assign n_11390 =  x_440 & ~n_11387;
assign n_11391 = ~n_11386 &  n_11390;
assign n_11392 =  n_10523 & ~n_11391;
assign n_11393 = ~n_11389 &  n_11392;
assign n_11394 = ~x_216 &  n_11346;
assign n_11395 =  x_216 & ~n_11346;
assign n_11396 = ~n_11394 & ~n_11395;
assign n_11397 = ~n_11350 & ~n_11354;
assign n_11398 =  n_11396 & ~n_11397;
assign n_11399 = ~n_11396 &  n_11397;
assign n_11400 = ~n_11398 & ~n_11399;
assign n_11401 = ~x_2680 & ~n_11400;
assign n_11402 =  x_2680 & ~n_11399;
assign n_11403 = ~n_11398 &  n_11402;
assign n_11404 =  n_10519 & ~n_11403;
assign n_11405 = ~n_11401 &  n_11404;
assign n_11406 = ~n_11393 & ~n_11405;
assign n_11407 =  n_11381 &  n_11406;
assign n_11408 =  x_1080 & ~n_11407;
assign n_11409 = ~x_1080 &  n_11407;
assign n_11410 = ~n_11408 & ~n_11409;
assign n_11411 = ~x_1687 &  n_11363;
assign n_11412 =  x_1687 & ~n_11363;
assign n_11413 = ~n_11411 & ~n_11412;
assign n_11414 = ~n_11367 & ~n_11371;
assign n_11415 =  n_11413 & ~n_11414;
assign n_11416 = ~n_11413 &  n_11414;
assign n_11417 = ~n_11415 & ~n_11416;
assign n_11418 = ~x_247 & ~n_11417;
assign n_11419 =  x_247 & ~n_11416;
assign n_11420 = ~n_11415 &  n_11419;
assign n_11421 =  n_10522 & ~n_11420;
assign n_11422 = ~n_11418 &  n_11421;
assign n_11423 =  x_1079 &  n_10525;
assign n_11424 =  x_855 & ~n_11377;
assign n_11425 = ~x_855 &  n_11377;
assign n_11426 =  n_10517 & ~n_11425;
assign n_11427 = ~n_11424 &  n_11426;
assign n_11428 = ~n_11423 & ~n_11427;
assign n_11429 = ~n_11422 &  n_11428;
assign n_11430 = ~x_2327 &  n_11382;
assign n_11431 =  x_2327 & ~n_11382;
assign n_11432 = ~n_11430 & ~n_11431;
assign n_11433 = ~n_11386 & ~n_11390;
assign n_11434 =  n_11432 & ~n_11433;
assign n_11435 = ~n_11432 &  n_11433;
assign n_11436 = ~n_11434 & ~n_11435;
assign n_11437 = ~x_439 & ~n_11436;
assign n_11438 =  x_439 & ~n_11435;
assign n_11439 = ~n_11434 &  n_11438;
assign n_11440 =  n_10523 & ~n_11439;
assign n_11441 = ~n_11437 &  n_11440;
assign n_11442 = ~x_215 &  n_11394;
assign n_11443 =  x_215 & ~n_11394;
assign n_11444 = ~n_11442 & ~n_11443;
assign n_11445 = ~n_11398 & ~n_11402;
assign n_11446 =  n_11444 & ~n_11445;
assign n_11447 = ~n_11444 &  n_11445;
assign n_11448 = ~n_11446 & ~n_11447;
assign n_11449 = ~x_2679 & ~n_11448;
assign n_11450 =  x_2679 & ~n_11447;
assign n_11451 = ~n_11446 &  n_11450;
assign n_11452 =  n_10519 & ~n_11451;
assign n_11453 = ~n_11449 &  n_11452;
assign n_11454 = ~n_11441 & ~n_11453;
assign n_11455 =  n_11429 &  n_11454;
assign n_11456 =  x_1079 & ~n_11455;
assign n_11457 = ~x_1079 &  n_11455;
assign n_11458 = ~n_11456 & ~n_11457;
assign n_11459 = ~x_1686 &  n_11411;
assign n_11460 =  x_1686 & ~n_11411;
assign n_11461 = ~n_11459 & ~n_11460;
assign n_11462 = ~n_11415 & ~n_11419;
assign n_11463 =  n_11461 & ~n_11462;
assign n_11464 = ~n_11461 &  n_11462;
assign n_11465 = ~n_11463 & ~n_11464;
assign n_11466 = ~x_246 & ~n_11465;
assign n_11467 =  x_246 & ~n_11464;
assign n_11468 = ~n_11463 &  n_11467;
assign n_11469 =  n_10522 & ~n_11468;
assign n_11470 = ~n_11466 &  n_11469;
assign n_11471 =  x_1078 &  n_10525;
assign n_11472 =  x_854 & ~n_11425;
assign n_11473 = ~x_854 &  n_11425;
assign n_11474 =  n_10517 & ~n_11473;
assign n_11475 = ~n_11472 &  n_11474;
assign n_11476 = ~n_11471 & ~n_11475;
assign n_11477 = ~n_11470 &  n_11476;
assign n_11478 = ~x_2326 &  n_11430;
assign n_11479 =  x_2326 & ~n_11430;
assign n_11480 = ~n_11478 & ~n_11479;
assign n_11481 = ~n_11434 & ~n_11438;
assign n_11482 =  n_11480 & ~n_11481;
assign n_11483 = ~n_11480 &  n_11481;
assign n_11484 = ~n_11482 & ~n_11483;
assign n_11485 = ~x_438 & ~n_11484;
assign n_11486 =  x_438 & ~n_11483;
assign n_11487 = ~n_11482 &  n_11486;
assign n_11488 =  n_10523 & ~n_11487;
assign n_11489 = ~n_11485 &  n_11488;
assign n_11490 = ~x_214 &  n_11442;
assign n_11491 =  x_214 & ~n_11442;
assign n_11492 = ~n_11490 & ~n_11491;
assign n_11493 = ~n_11446 & ~n_11450;
assign n_11494 =  n_11492 & ~n_11493;
assign n_11495 = ~n_11492 &  n_11493;
assign n_11496 = ~n_11494 & ~n_11495;
assign n_11497 = ~x_2678 & ~n_11496;
assign n_11498 =  x_2678 & ~n_11495;
assign n_11499 = ~n_11494 &  n_11498;
assign n_11500 =  n_10519 & ~n_11499;
assign n_11501 = ~n_11497 &  n_11500;
assign n_11502 = ~n_11489 & ~n_11501;
assign n_11503 =  n_11477 &  n_11502;
assign n_11504 =  x_1078 & ~n_11503;
assign n_11505 = ~x_1078 &  n_11503;
assign n_11506 = ~n_11504 & ~n_11505;
assign n_11507 = ~x_1685 &  n_11459;
assign n_11508 =  x_1685 & ~n_11459;
assign n_11509 = ~n_11507 & ~n_11508;
assign n_11510 = ~n_11463 & ~n_11467;
assign n_11511 =  n_11509 & ~n_11510;
assign n_11512 = ~n_11509 &  n_11510;
assign n_11513 = ~n_11511 & ~n_11512;
assign n_11514 = ~x_245 & ~n_11513;
assign n_11515 =  x_245 & ~n_11512;
assign n_11516 = ~n_11511 &  n_11515;
assign n_11517 =  n_10522 & ~n_11516;
assign n_11518 = ~n_11514 &  n_11517;
assign n_11519 =  x_1077 &  n_10525;
assign n_11520 =  x_853 & ~n_11473;
assign n_11521 = ~x_853 &  n_11473;
assign n_11522 =  n_10517 & ~n_11521;
assign n_11523 = ~n_11520 &  n_11522;
assign n_11524 = ~n_11519 & ~n_11523;
assign n_11525 = ~n_11518 &  n_11524;
assign n_11526 = ~x_2325 &  n_11478;
assign n_11527 =  x_2325 & ~n_11478;
assign n_11528 = ~n_11526 & ~n_11527;
assign n_11529 = ~n_11482 & ~n_11486;
assign n_11530 =  n_11528 & ~n_11529;
assign n_11531 = ~n_11528 &  n_11529;
assign n_11532 = ~n_11530 & ~n_11531;
assign n_11533 = ~x_437 & ~n_11532;
assign n_11534 =  x_437 & ~n_11531;
assign n_11535 = ~n_11530 &  n_11534;
assign n_11536 =  n_10523 & ~n_11535;
assign n_11537 = ~n_11533 &  n_11536;
assign n_11538 = ~x_213 &  n_11490;
assign n_11539 =  x_213 & ~n_11490;
assign n_11540 = ~n_11538 & ~n_11539;
assign n_11541 = ~n_11494 & ~n_11498;
assign n_11542 =  n_11540 & ~n_11541;
assign n_11543 = ~n_11540 &  n_11541;
assign n_11544 = ~n_11542 & ~n_11543;
assign n_11545 = ~x_2677 & ~n_11544;
assign n_11546 =  x_2677 & ~n_11543;
assign n_11547 = ~n_11542 &  n_11546;
assign n_11548 =  n_10519 & ~n_11547;
assign n_11549 = ~n_11545 &  n_11548;
assign n_11550 = ~n_11537 & ~n_11549;
assign n_11551 =  n_11525 &  n_11550;
assign n_11552 =  x_1077 & ~n_11551;
assign n_11553 = ~x_1077 &  n_11551;
assign n_11554 = ~n_11552 & ~n_11553;
assign n_11555 = ~x_1684 &  n_11507;
assign n_11556 =  x_1684 & ~n_11507;
assign n_11557 = ~n_11555 & ~n_11556;
assign n_11558 = ~n_11511 & ~n_11515;
assign n_11559 =  n_11557 & ~n_11558;
assign n_11560 = ~n_11557 &  n_11558;
assign n_11561 = ~n_11559 & ~n_11560;
assign n_11562 = ~x_244 & ~n_11561;
assign n_11563 =  x_244 & ~n_11560;
assign n_11564 = ~n_11559 &  n_11563;
assign n_11565 =  n_10522 & ~n_11564;
assign n_11566 = ~n_11562 &  n_11565;
assign n_11567 =  x_1076 &  n_10525;
assign n_11568 =  x_852 & ~n_11521;
assign n_11569 = ~x_852 &  n_11521;
assign n_11570 =  n_10517 & ~n_11569;
assign n_11571 = ~n_11568 &  n_11570;
assign n_11572 = ~n_11567 & ~n_11571;
assign n_11573 = ~n_11566 &  n_11572;
assign n_11574 = ~x_2324 &  n_11526;
assign n_11575 =  x_2324 & ~n_11526;
assign n_11576 = ~n_11574 & ~n_11575;
assign n_11577 = ~n_11530 & ~n_11534;
assign n_11578 =  n_11576 & ~n_11577;
assign n_11579 = ~n_11576 &  n_11577;
assign n_11580 = ~n_11578 & ~n_11579;
assign n_11581 = ~x_436 & ~n_11580;
assign n_11582 =  x_436 & ~n_11579;
assign n_11583 = ~n_11578 &  n_11582;
assign n_11584 =  n_10523 & ~n_11583;
assign n_11585 = ~n_11581 &  n_11584;
assign n_11586 = ~x_212 &  n_11538;
assign n_11587 =  x_212 & ~n_11538;
assign n_11588 = ~n_11586 & ~n_11587;
assign n_11589 = ~n_11542 & ~n_11546;
assign n_11590 =  n_11588 & ~n_11589;
assign n_11591 = ~n_11588 &  n_11589;
assign n_11592 = ~n_11590 & ~n_11591;
assign n_11593 = ~x_2676 & ~n_11592;
assign n_11594 =  x_2676 & ~n_11591;
assign n_11595 = ~n_11590 &  n_11594;
assign n_11596 =  n_10519 & ~n_11595;
assign n_11597 = ~n_11593 &  n_11596;
assign n_11598 = ~n_11585 & ~n_11597;
assign n_11599 =  n_11573 &  n_11598;
assign n_11600 =  x_1076 & ~n_11599;
assign n_11601 = ~x_1076 &  n_11599;
assign n_11602 = ~n_11600 & ~n_11601;
assign n_11603 = ~x_1683 &  n_11555;
assign n_11604 =  x_1683 & ~n_11555;
assign n_11605 = ~n_11603 & ~n_11604;
assign n_11606 = ~n_11559 & ~n_11563;
assign n_11607 =  n_11605 & ~n_11606;
assign n_11608 = ~n_11605 &  n_11606;
assign n_11609 = ~n_11607 & ~n_11608;
assign n_11610 = ~x_243 & ~n_11609;
assign n_11611 =  x_243 & ~n_11608;
assign n_11612 = ~n_11607 &  n_11611;
assign n_11613 =  n_10522 & ~n_11612;
assign n_11614 = ~n_11610 &  n_11613;
assign n_11615 =  x_1075 &  n_10525;
assign n_11616 =  x_851 & ~n_11569;
assign n_11617 = ~x_851 &  n_11569;
assign n_11618 =  n_10517 & ~n_11617;
assign n_11619 = ~n_11616 &  n_11618;
assign n_11620 = ~n_11615 & ~n_11619;
assign n_11621 = ~n_11614 &  n_11620;
assign n_11622 = ~x_2323 &  n_11574;
assign n_11623 =  x_2323 & ~n_11574;
assign n_11624 = ~n_11622 & ~n_11623;
assign n_11625 = ~n_11578 & ~n_11582;
assign n_11626 =  n_11624 & ~n_11625;
assign n_11627 = ~n_11624 &  n_11625;
assign n_11628 = ~n_11626 & ~n_11627;
assign n_11629 = ~x_435 & ~n_11628;
assign n_11630 =  x_435 & ~n_11627;
assign n_11631 = ~n_11626 &  n_11630;
assign n_11632 =  n_10523 & ~n_11631;
assign n_11633 = ~n_11629 &  n_11632;
assign n_11634 = ~x_211 &  n_11586;
assign n_11635 =  x_211 & ~n_11586;
assign n_11636 = ~n_11634 & ~n_11635;
assign n_11637 = ~n_11590 & ~n_11594;
assign n_11638 =  n_11636 & ~n_11637;
assign n_11639 = ~n_11636 &  n_11637;
assign n_11640 = ~n_11638 & ~n_11639;
assign n_11641 = ~x_2675 & ~n_11640;
assign n_11642 =  x_2675 & ~n_11639;
assign n_11643 = ~n_11638 &  n_11642;
assign n_11644 =  n_10519 & ~n_11643;
assign n_11645 = ~n_11641 &  n_11644;
assign n_11646 = ~n_11633 & ~n_11645;
assign n_11647 =  n_11621 &  n_11646;
assign n_11648 =  x_1075 & ~n_11647;
assign n_11649 = ~x_1075 &  n_11647;
assign n_11650 = ~n_11648 & ~n_11649;
assign n_11651 = ~x_1682 &  n_11603;
assign n_11652 =  x_1682 & ~n_11603;
assign n_11653 = ~n_11651 & ~n_11652;
assign n_11654 = ~n_11607 & ~n_11611;
assign n_11655 =  n_11653 & ~n_11654;
assign n_11656 = ~n_11653 &  n_11654;
assign n_11657 = ~n_11655 & ~n_11656;
assign n_11658 = ~x_242 & ~n_11657;
assign n_11659 =  x_242 & ~n_11656;
assign n_11660 = ~n_11655 &  n_11659;
assign n_11661 =  n_10522 & ~n_11660;
assign n_11662 = ~n_11658 &  n_11661;
assign n_11663 =  x_1074 &  n_10525;
assign n_11664 =  x_850 & ~n_11617;
assign n_11665 = ~x_850 &  n_11617;
assign n_11666 =  n_10517 & ~n_11665;
assign n_11667 = ~n_11664 &  n_11666;
assign n_11668 = ~n_11663 & ~n_11667;
assign n_11669 = ~n_11662 &  n_11668;
assign n_11670 = ~x_2322 &  n_11622;
assign n_11671 =  x_2322 & ~n_11622;
assign n_11672 = ~n_11670 & ~n_11671;
assign n_11673 = ~n_11626 & ~n_11630;
assign n_11674 =  n_11672 & ~n_11673;
assign n_11675 = ~n_11672 &  n_11673;
assign n_11676 = ~n_11674 & ~n_11675;
assign n_11677 = ~x_434 & ~n_11676;
assign n_11678 =  x_434 & ~n_11675;
assign n_11679 = ~n_11674 &  n_11678;
assign n_11680 =  n_10523 & ~n_11679;
assign n_11681 = ~n_11677 &  n_11680;
assign n_11682 = ~x_210 &  n_11634;
assign n_11683 =  x_210 & ~n_11634;
assign n_11684 = ~n_11682 & ~n_11683;
assign n_11685 = ~n_11638 & ~n_11642;
assign n_11686 =  n_11684 & ~n_11685;
assign n_11687 = ~n_11684 &  n_11685;
assign n_11688 = ~n_11686 & ~n_11687;
assign n_11689 = ~x_2674 & ~n_11688;
assign n_11690 =  x_2674 & ~n_11687;
assign n_11691 = ~n_11686 &  n_11690;
assign n_11692 =  n_10519 & ~n_11691;
assign n_11693 = ~n_11689 &  n_11692;
assign n_11694 = ~n_11681 & ~n_11693;
assign n_11695 =  n_11669 &  n_11694;
assign n_11696 =  x_1074 & ~n_11695;
assign n_11697 = ~x_1074 &  n_11695;
assign n_11698 = ~n_11696 & ~n_11697;
assign n_11699 = ~x_1681 &  n_11651;
assign n_11700 =  x_1681 & ~n_11651;
assign n_11701 = ~n_11699 & ~n_11700;
assign n_11702 = ~n_11655 & ~n_11659;
assign n_11703 =  n_11701 & ~n_11702;
assign n_11704 = ~n_11701 &  n_11702;
assign n_11705 = ~n_11703 & ~n_11704;
assign n_11706 = ~x_241 & ~n_11705;
assign n_11707 =  x_241 & ~n_11704;
assign n_11708 = ~n_11703 &  n_11707;
assign n_11709 =  n_10522 & ~n_11708;
assign n_11710 = ~n_11706 &  n_11709;
assign n_11711 =  x_1073 &  n_10525;
assign n_11712 =  x_849 & ~n_11665;
assign n_11713 = ~x_849 &  n_11665;
assign n_11714 =  n_10517 & ~n_11713;
assign n_11715 = ~n_11712 &  n_11714;
assign n_11716 = ~n_11711 & ~n_11715;
assign n_11717 = ~n_11710 &  n_11716;
assign n_11718 = ~x_2321 &  n_11670;
assign n_11719 =  x_2321 & ~n_11670;
assign n_11720 = ~n_11718 & ~n_11719;
assign n_11721 = ~n_11674 & ~n_11678;
assign n_11722 =  n_11720 & ~n_11721;
assign n_11723 = ~n_11720 &  n_11721;
assign n_11724 = ~n_11722 & ~n_11723;
assign n_11725 = ~x_433 & ~n_11724;
assign n_11726 =  x_433 & ~n_11723;
assign n_11727 = ~n_11722 &  n_11726;
assign n_11728 =  n_10523 & ~n_11727;
assign n_11729 = ~n_11725 &  n_11728;
assign n_11730 = ~x_209 &  n_11682;
assign n_11731 =  x_209 & ~n_11682;
assign n_11732 = ~n_11730 & ~n_11731;
assign n_11733 = ~n_11686 & ~n_11690;
assign n_11734 =  n_11732 & ~n_11733;
assign n_11735 = ~n_11732 &  n_11733;
assign n_11736 = ~n_11734 & ~n_11735;
assign n_11737 = ~x_2673 & ~n_11736;
assign n_11738 =  x_2673 & ~n_11735;
assign n_11739 = ~n_11734 &  n_11738;
assign n_11740 =  n_10519 & ~n_11739;
assign n_11741 = ~n_11737 &  n_11740;
assign n_11742 = ~n_11729 & ~n_11741;
assign n_11743 =  n_11717 &  n_11742;
assign n_11744 =  x_1073 & ~n_11743;
assign n_11745 = ~x_1073 &  n_11743;
assign n_11746 = ~n_11744 & ~n_11745;
assign n_11747 = ~x_1680 &  n_11699;
assign n_11748 =  x_1680 & ~n_11699;
assign n_11749 = ~n_11747 & ~n_11748;
assign n_11750 = ~n_11703 & ~n_11707;
assign n_11751 =  n_11749 & ~n_11750;
assign n_11752 = ~n_11749 &  n_11750;
assign n_11753 = ~n_11751 & ~n_11752;
assign n_11754 = ~x_240 & ~n_11753;
assign n_11755 =  x_240 & ~n_11752;
assign n_11756 = ~n_11751 &  n_11755;
assign n_11757 =  n_10522 & ~n_11756;
assign n_11758 = ~n_11754 &  n_11757;
assign n_11759 =  x_1072 &  n_10525;
assign n_11760 =  x_848 & ~n_11713;
assign n_11761 = ~x_848 &  n_11713;
assign n_11762 =  n_10517 & ~n_11761;
assign n_11763 = ~n_11760 &  n_11762;
assign n_11764 = ~n_11759 & ~n_11763;
assign n_11765 = ~n_11758 &  n_11764;
assign n_11766 = ~x_2320 &  n_11718;
assign n_11767 =  x_2320 & ~n_11718;
assign n_11768 = ~n_11766 & ~n_11767;
assign n_11769 = ~n_11722 & ~n_11726;
assign n_11770 =  n_11768 & ~n_11769;
assign n_11771 = ~n_11768 &  n_11769;
assign n_11772 = ~n_11770 & ~n_11771;
assign n_11773 = ~x_432 & ~n_11772;
assign n_11774 =  x_432 & ~n_11771;
assign n_11775 = ~n_11770 &  n_11774;
assign n_11776 =  n_10523 & ~n_11775;
assign n_11777 = ~n_11773 &  n_11776;
assign n_11778 = ~x_208 &  n_11730;
assign n_11779 =  x_208 & ~n_11730;
assign n_11780 = ~n_11778 & ~n_11779;
assign n_11781 = ~n_11734 & ~n_11738;
assign n_11782 =  n_11780 & ~n_11781;
assign n_11783 = ~n_11780 &  n_11781;
assign n_11784 = ~n_11782 & ~n_11783;
assign n_11785 = ~x_2672 & ~n_11784;
assign n_11786 =  x_2672 & ~n_11783;
assign n_11787 = ~n_11782 &  n_11786;
assign n_11788 =  n_10519 & ~n_11787;
assign n_11789 = ~n_11785 &  n_11788;
assign n_11790 = ~n_11777 & ~n_11789;
assign n_11791 =  n_11765 &  n_11790;
assign n_11792 =  x_1072 & ~n_11791;
assign n_11793 = ~x_1072 &  n_11791;
assign n_11794 = ~n_11792 & ~n_11793;
assign n_11795 = ~x_1679 &  n_11747;
assign n_11796 =  x_1679 & ~n_11747;
assign n_11797 = ~n_11795 & ~n_11796;
assign n_11798 = ~n_11751 & ~n_11755;
assign n_11799 =  n_11797 & ~n_11798;
assign n_11800 = ~n_11797 &  n_11798;
assign n_11801 = ~n_11799 & ~n_11800;
assign n_11802 = ~x_239 & ~n_11801;
assign n_11803 =  x_239 & ~n_11800;
assign n_11804 = ~n_11799 &  n_11803;
assign n_11805 =  n_10522 & ~n_11804;
assign n_11806 = ~n_11802 &  n_11805;
assign n_11807 =  x_1071 &  n_10525;
assign n_11808 =  x_847 & ~n_11761;
assign n_11809 = ~x_847 &  n_11761;
assign n_11810 =  n_10517 & ~n_11809;
assign n_11811 = ~n_11808 &  n_11810;
assign n_11812 = ~n_11807 & ~n_11811;
assign n_11813 = ~n_11806 &  n_11812;
assign n_11814 = ~x_2319 &  n_11766;
assign n_11815 =  x_2319 & ~n_11766;
assign n_11816 = ~n_11814 & ~n_11815;
assign n_11817 = ~n_11770 & ~n_11774;
assign n_11818 =  n_11816 & ~n_11817;
assign n_11819 = ~n_11816 &  n_11817;
assign n_11820 = ~n_11818 & ~n_11819;
assign n_11821 = ~x_431 & ~n_11820;
assign n_11822 =  x_431 & ~n_11819;
assign n_11823 = ~n_11818 &  n_11822;
assign n_11824 =  n_10523 & ~n_11823;
assign n_11825 = ~n_11821 &  n_11824;
assign n_11826 = ~x_207 &  n_11778;
assign n_11827 =  x_207 & ~n_11778;
assign n_11828 = ~n_11826 & ~n_11827;
assign n_11829 = ~n_11782 & ~n_11786;
assign n_11830 =  n_11828 & ~n_11829;
assign n_11831 = ~n_11828 &  n_11829;
assign n_11832 = ~n_11830 & ~n_11831;
assign n_11833 = ~x_2671 & ~n_11832;
assign n_11834 =  x_2671 & ~n_11831;
assign n_11835 = ~n_11830 &  n_11834;
assign n_11836 =  n_10519 & ~n_11835;
assign n_11837 = ~n_11833 &  n_11836;
assign n_11838 = ~n_11825 & ~n_11837;
assign n_11839 =  n_11813 &  n_11838;
assign n_11840 =  x_1071 & ~n_11839;
assign n_11841 = ~x_1071 &  n_11839;
assign n_11842 = ~n_11840 & ~n_11841;
assign n_11843 = ~x_1678 &  n_11795;
assign n_11844 =  x_1678 & ~n_11795;
assign n_11845 = ~n_11843 & ~n_11844;
assign n_11846 = ~n_11799 & ~n_11803;
assign n_11847 =  n_11845 & ~n_11846;
assign n_11848 = ~n_11845 &  n_11846;
assign n_11849 = ~n_11847 & ~n_11848;
assign n_11850 = ~x_238 & ~n_11849;
assign n_11851 =  x_238 & ~n_11848;
assign n_11852 = ~n_11847 &  n_11851;
assign n_11853 =  n_10522 & ~n_11852;
assign n_11854 = ~n_11850 &  n_11853;
assign n_11855 =  x_1070 &  n_10525;
assign n_11856 =  x_846 & ~n_11809;
assign n_11857 = ~x_846 &  n_11809;
assign n_11858 =  n_10517 & ~n_11857;
assign n_11859 = ~n_11856 &  n_11858;
assign n_11860 = ~n_11855 & ~n_11859;
assign n_11861 = ~n_11854 &  n_11860;
assign n_11862 = ~x_2318 &  n_11814;
assign n_11863 =  x_2318 & ~n_11814;
assign n_11864 = ~n_11862 & ~n_11863;
assign n_11865 = ~n_11818 & ~n_11822;
assign n_11866 =  n_11864 & ~n_11865;
assign n_11867 = ~n_11864 &  n_11865;
assign n_11868 = ~n_11866 & ~n_11867;
assign n_11869 = ~x_430 & ~n_11868;
assign n_11870 =  x_430 & ~n_11867;
assign n_11871 = ~n_11866 &  n_11870;
assign n_11872 =  n_10523 & ~n_11871;
assign n_11873 = ~n_11869 &  n_11872;
assign n_11874 = ~x_206 &  n_11826;
assign n_11875 =  x_206 & ~n_11826;
assign n_11876 = ~n_11874 & ~n_11875;
assign n_11877 = ~n_11830 & ~n_11834;
assign n_11878 =  n_11876 & ~n_11877;
assign n_11879 = ~n_11876 &  n_11877;
assign n_11880 = ~n_11878 & ~n_11879;
assign n_11881 = ~x_2670 & ~n_11880;
assign n_11882 =  x_2670 & ~n_11879;
assign n_11883 = ~n_11878 &  n_11882;
assign n_11884 =  n_10519 & ~n_11883;
assign n_11885 = ~n_11881 &  n_11884;
assign n_11886 = ~n_11873 & ~n_11885;
assign n_11887 =  n_11861 &  n_11886;
assign n_11888 =  x_1070 & ~n_11887;
assign n_11889 = ~x_1070 &  n_11887;
assign n_11890 = ~n_11888 & ~n_11889;
assign n_11891 = ~x_1677 &  n_11843;
assign n_11892 =  x_1677 & ~n_11843;
assign n_11893 = ~n_11891 & ~n_11892;
assign n_11894 = ~n_11847 & ~n_11851;
assign n_11895 =  n_11893 & ~n_11894;
assign n_11896 = ~n_11893 &  n_11894;
assign n_11897 = ~n_11895 & ~n_11896;
assign n_11898 = ~x_237 & ~n_11897;
assign n_11899 =  x_237 & ~n_11896;
assign n_11900 = ~n_11895 &  n_11899;
assign n_11901 =  n_10522 & ~n_11900;
assign n_11902 = ~n_11898 &  n_11901;
assign n_11903 =  x_1069 &  n_10525;
assign n_11904 =  x_845 & ~n_11857;
assign n_11905 = ~x_845 &  n_11857;
assign n_11906 =  n_10517 & ~n_11905;
assign n_11907 = ~n_11904 &  n_11906;
assign n_11908 = ~n_11903 & ~n_11907;
assign n_11909 = ~n_11902 &  n_11908;
assign n_11910 = ~x_2317 &  n_11862;
assign n_11911 =  x_2317 & ~n_11862;
assign n_11912 = ~n_11910 & ~n_11911;
assign n_11913 = ~n_11866 & ~n_11870;
assign n_11914 =  n_11912 & ~n_11913;
assign n_11915 = ~n_11912 &  n_11913;
assign n_11916 = ~n_11914 & ~n_11915;
assign n_11917 = ~x_429 & ~n_11916;
assign n_11918 =  x_429 & ~n_11915;
assign n_11919 = ~n_11914 &  n_11918;
assign n_11920 =  n_10523 & ~n_11919;
assign n_11921 = ~n_11917 &  n_11920;
assign n_11922 = ~x_205 &  n_11874;
assign n_11923 =  x_205 & ~n_11874;
assign n_11924 = ~n_11922 & ~n_11923;
assign n_11925 = ~n_11878 & ~n_11882;
assign n_11926 =  n_11924 & ~n_11925;
assign n_11927 = ~n_11924 &  n_11925;
assign n_11928 = ~n_11926 & ~n_11927;
assign n_11929 = ~x_2669 & ~n_11928;
assign n_11930 =  x_2669 & ~n_11927;
assign n_11931 = ~n_11926 &  n_11930;
assign n_11932 =  n_10519 & ~n_11931;
assign n_11933 = ~n_11929 &  n_11932;
assign n_11934 = ~n_11921 & ~n_11933;
assign n_11935 =  n_11909 &  n_11934;
assign n_11936 =  x_1069 & ~n_11935;
assign n_11937 = ~x_1069 &  n_11935;
assign n_11938 = ~n_11936 & ~n_11937;
assign n_11939 = ~x_1676 &  n_11891;
assign n_11940 =  x_1676 & ~n_11891;
assign n_11941 = ~n_11939 & ~n_11940;
assign n_11942 = ~n_11895 & ~n_11899;
assign n_11943 =  n_11941 & ~n_11942;
assign n_11944 = ~n_11941 &  n_11942;
assign n_11945 = ~n_11943 & ~n_11944;
assign n_11946 = ~x_236 & ~n_11945;
assign n_11947 =  x_236 & ~n_11944;
assign n_11948 = ~n_11943 &  n_11947;
assign n_11949 =  n_10522 & ~n_11948;
assign n_11950 = ~n_11946 &  n_11949;
assign n_11951 =  x_1068 &  n_10525;
assign n_11952 =  x_844 & ~n_11905;
assign n_11953 = ~x_844 &  n_11905;
assign n_11954 =  n_10517 & ~n_11953;
assign n_11955 = ~n_11952 &  n_11954;
assign n_11956 = ~n_11951 & ~n_11955;
assign n_11957 = ~n_11950 &  n_11956;
assign n_11958 = ~x_2316 &  n_11910;
assign n_11959 =  x_2316 & ~n_11910;
assign n_11960 = ~n_11958 & ~n_11959;
assign n_11961 = ~n_11914 & ~n_11918;
assign n_11962 =  n_11960 & ~n_11961;
assign n_11963 = ~n_11960 &  n_11961;
assign n_11964 = ~n_11962 & ~n_11963;
assign n_11965 = ~x_428 & ~n_11964;
assign n_11966 =  x_428 & ~n_11963;
assign n_11967 = ~n_11962 &  n_11966;
assign n_11968 =  n_10523 & ~n_11967;
assign n_11969 = ~n_11965 &  n_11968;
assign n_11970 = ~x_204 &  n_11922;
assign n_11971 =  x_204 & ~n_11922;
assign n_11972 = ~n_11970 & ~n_11971;
assign n_11973 = ~n_11926 & ~n_11930;
assign n_11974 =  n_11972 & ~n_11973;
assign n_11975 = ~n_11972 &  n_11973;
assign n_11976 = ~n_11974 & ~n_11975;
assign n_11977 = ~x_2668 & ~n_11976;
assign n_11978 =  x_2668 & ~n_11975;
assign n_11979 = ~n_11974 &  n_11978;
assign n_11980 =  n_10519 & ~n_11979;
assign n_11981 = ~n_11977 &  n_11980;
assign n_11982 = ~n_11969 & ~n_11981;
assign n_11983 =  n_11957 &  n_11982;
assign n_11984 =  x_1068 & ~n_11983;
assign n_11985 = ~x_1068 &  n_11983;
assign n_11986 = ~n_11984 & ~n_11985;
assign n_11987 = ~n_11962 & ~n_11966;
assign n_11988 =  x_427 & ~x_2315;
assign n_11989 = ~x_427 &  x_2315;
assign n_11990 = ~n_11988 & ~n_11989;
assign n_11991 =  n_11958 &  n_11990;
assign n_11992 = ~n_11958 & ~n_11990;
assign n_11993 = ~n_11991 & ~n_11992;
assign n_11994 =  n_11987 & ~n_11993;
assign n_11995 = ~n_11987 &  n_11993;
assign n_11996 =  n_10523 & ~n_11995;
assign n_11997 = ~n_11994 &  n_11996;
assign n_11998 =  x_1067 &  n_10525;
assign n_11999 = ~x_843 &  n_11953;
assign n_12000 =  x_843 & ~n_11953;
assign n_12001 =  n_10517 & ~n_12000;
assign n_12002 = ~n_11999 &  n_12001;
assign n_12003 = ~n_11998 & ~n_12002;
assign n_12004 = ~n_11997 &  n_12003;
assign n_12005 = ~n_11974 & ~n_11978;
assign n_12006 =  x_203 & ~x_2667;
assign n_12007 = ~x_203 &  x_2667;
assign n_12008 = ~n_12006 & ~n_12007;
assign n_12009 =  n_11970 &  n_12008;
assign n_12010 = ~n_11970 & ~n_12008;
assign n_12011 = ~n_12009 & ~n_12010;
assign n_12012 =  n_12005 & ~n_12011;
assign n_12013 = ~n_12005 &  n_12011;
assign n_12014 =  n_10519 & ~n_12013;
assign n_12015 = ~n_12012 &  n_12014;
assign n_12016 = ~n_11943 & ~n_11947;
assign n_12017 =  x_235 & ~x_1675;
assign n_12018 = ~x_235 &  x_1675;
assign n_12019 = ~n_12017 & ~n_12018;
assign n_12020 =  n_11939 &  n_12019;
assign n_12021 = ~n_11939 & ~n_12019;
assign n_12022 = ~n_12020 & ~n_12021;
assign n_12023 =  n_12016 & ~n_12022;
assign n_12024 = ~n_12016 &  n_12022;
assign n_12025 =  n_10522 & ~n_12024;
assign n_12026 = ~n_12023 &  n_12025;
assign n_12027 = ~n_12015 & ~n_12026;
assign n_12028 =  n_12004 &  n_12027;
assign n_12029 =  x_1067 & ~n_12028;
assign n_12030 = ~x_1067 &  n_12028;
assign n_12031 = ~n_12029 & ~n_12030;
assign n_12032 =  n_10319 &  n_1903;
assign n_12033 =  n_586 &  n_12032;
assign n_12034 =  x_1066 & ~n_12033;
assign n_12035 =  x_426 &  n_12033;
assign n_12036 = ~n_12034 & ~n_12035;
assign n_12037 =  x_1066 & ~n_12036;
assign n_12038 = ~x_1066 &  n_12036;
assign n_12039 = ~n_12037 & ~n_12038;
assign n_12040 =  x_1065 & ~n_12033;
assign n_12041 =  x_425 &  n_12033;
assign n_12042 = ~n_12040 & ~n_12041;
assign n_12043 =  x_1065 & ~n_12042;
assign n_12044 = ~x_1065 &  n_12042;
assign n_12045 = ~n_12043 & ~n_12044;
assign n_12046 =  x_1064 & ~n_12033;
assign n_12047 =  x_424 &  n_12033;
assign n_12048 = ~n_12046 & ~n_12047;
assign n_12049 =  x_1064 & ~n_12048;
assign n_12050 = ~x_1064 &  n_12048;
assign n_12051 = ~n_12049 & ~n_12050;
assign n_12052 =  x_1063 & ~n_12033;
assign n_12053 =  x_423 &  n_12033;
assign n_12054 = ~n_12052 & ~n_12053;
assign n_12055 =  x_1063 & ~n_12054;
assign n_12056 = ~x_1063 &  n_12054;
assign n_12057 = ~n_12055 & ~n_12056;
assign n_12058 =  x_1062 & ~n_12033;
assign n_12059 =  x_422 &  n_12033;
assign n_12060 = ~n_12058 & ~n_12059;
assign n_12061 =  x_1062 & ~n_12060;
assign n_12062 = ~x_1062 &  n_12060;
assign n_12063 = ~n_12061 & ~n_12062;
assign n_12064 =  x_1061 & ~n_12033;
assign n_12065 =  x_421 &  n_12033;
assign n_12066 = ~n_12064 & ~n_12065;
assign n_12067 =  x_1061 & ~n_12066;
assign n_12068 = ~x_1061 &  n_12066;
assign n_12069 = ~n_12067 & ~n_12068;
assign n_12070 =  x_1060 & ~n_12033;
assign n_12071 =  x_420 &  n_12033;
assign n_12072 = ~n_12070 & ~n_12071;
assign n_12073 =  x_1060 & ~n_12072;
assign n_12074 = ~x_1060 &  n_12072;
assign n_12075 = ~n_12073 & ~n_12074;
assign n_12076 =  x_1059 & ~n_12033;
assign n_12077 =  x_419 &  n_12033;
assign n_12078 = ~n_12076 & ~n_12077;
assign n_12079 =  x_1059 & ~n_12078;
assign n_12080 = ~x_1059 &  n_12078;
assign n_12081 = ~n_12079 & ~n_12080;
assign n_12082 =  x_1058 & ~n_12033;
assign n_12083 =  x_418 &  n_12033;
assign n_12084 = ~n_12082 & ~n_12083;
assign n_12085 =  x_1058 & ~n_12084;
assign n_12086 = ~x_1058 &  n_12084;
assign n_12087 = ~n_12085 & ~n_12086;
assign n_12088 =  x_1057 & ~n_12033;
assign n_12089 =  x_417 &  n_12033;
assign n_12090 = ~n_12088 & ~n_12089;
assign n_12091 =  x_1057 & ~n_12090;
assign n_12092 = ~x_1057 &  n_12090;
assign n_12093 = ~n_12091 & ~n_12092;
assign n_12094 =  x_1056 & ~n_12033;
assign n_12095 =  x_416 &  n_12033;
assign n_12096 = ~n_12094 & ~n_12095;
assign n_12097 =  x_1056 & ~n_12096;
assign n_12098 = ~x_1056 &  n_12096;
assign n_12099 = ~n_12097 & ~n_12098;
assign n_12100 =  x_1055 & ~n_12033;
assign n_12101 =  x_415 &  n_12033;
assign n_12102 = ~n_12100 & ~n_12101;
assign n_12103 =  x_1055 & ~n_12102;
assign n_12104 = ~x_1055 &  n_12102;
assign n_12105 = ~n_12103 & ~n_12104;
assign n_12106 =  x_1054 & ~n_12033;
assign n_12107 =  x_414 &  n_12033;
assign n_12108 = ~n_12106 & ~n_12107;
assign n_12109 =  x_1054 & ~n_12108;
assign n_12110 = ~x_1054 &  n_12108;
assign n_12111 = ~n_12109 & ~n_12110;
assign n_12112 =  x_1053 & ~n_12033;
assign n_12113 =  x_413 &  n_12033;
assign n_12114 = ~n_12112 & ~n_12113;
assign n_12115 =  x_1053 & ~n_12114;
assign n_12116 = ~x_1053 &  n_12114;
assign n_12117 = ~n_12115 & ~n_12116;
assign n_12118 =  x_1052 & ~n_12033;
assign n_12119 =  x_412 &  n_12033;
assign n_12120 = ~n_12118 & ~n_12119;
assign n_12121 =  x_1052 & ~n_12120;
assign n_12122 = ~x_1052 &  n_12120;
assign n_12123 = ~n_12121 & ~n_12122;
assign n_12124 =  x_1051 & ~n_12033;
assign n_12125 =  x_411 &  n_12033;
assign n_12126 = ~n_12124 & ~n_12125;
assign n_12127 =  x_1051 & ~n_12126;
assign n_12128 = ~x_1051 &  n_12126;
assign n_12129 = ~n_12127 & ~n_12128;
assign n_12130 =  x_1050 & ~n_12033;
assign n_12131 =  x_410 &  n_12033;
assign n_12132 = ~n_12130 & ~n_12131;
assign n_12133 =  x_1050 & ~n_12132;
assign n_12134 = ~x_1050 &  n_12132;
assign n_12135 = ~n_12133 & ~n_12134;
assign n_12136 =  x_1049 & ~n_12033;
assign n_12137 =  x_409 &  n_12033;
assign n_12138 = ~n_12136 & ~n_12137;
assign n_12139 =  x_1049 & ~n_12138;
assign n_12140 = ~x_1049 &  n_12138;
assign n_12141 = ~n_12139 & ~n_12140;
assign n_12142 =  x_1048 & ~n_12033;
assign n_12143 =  x_408 &  n_12033;
assign n_12144 = ~n_12142 & ~n_12143;
assign n_12145 =  x_1048 & ~n_12144;
assign n_12146 = ~x_1048 &  n_12144;
assign n_12147 = ~n_12145 & ~n_12146;
assign n_12148 =  x_1047 & ~n_12033;
assign n_12149 =  x_407 &  n_12033;
assign n_12150 = ~n_12148 & ~n_12149;
assign n_12151 =  x_1047 & ~n_12150;
assign n_12152 = ~x_1047 &  n_12150;
assign n_12153 = ~n_12151 & ~n_12152;
assign n_12154 =  x_1046 & ~n_12033;
assign n_12155 =  x_406 &  n_12033;
assign n_12156 = ~n_12154 & ~n_12155;
assign n_12157 =  x_1046 & ~n_12156;
assign n_12158 = ~x_1046 &  n_12156;
assign n_12159 = ~n_12157 & ~n_12158;
assign n_12160 =  x_1045 & ~n_12033;
assign n_12161 =  x_405 &  n_12033;
assign n_12162 = ~n_12160 & ~n_12161;
assign n_12163 =  x_1045 & ~n_12162;
assign n_12164 = ~x_1045 &  n_12162;
assign n_12165 = ~n_12163 & ~n_12164;
assign n_12166 =  x_1044 & ~n_12033;
assign n_12167 =  x_404 &  n_12033;
assign n_12168 = ~n_12166 & ~n_12167;
assign n_12169 =  x_1044 & ~n_12168;
assign n_12170 = ~x_1044 &  n_12168;
assign n_12171 = ~n_12169 & ~n_12170;
assign n_12172 =  x_1043 & ~n_12033;
assign n_12173 =  x_403 &  n_12033;
assign n_12174 = ~n_12172 & ~n_12173;
assign n_12175 =  x_1043 & ~n_12174;
assign n_12176 = ~x_1043 &  n_12174;
assign n_12177 = ~n_12175 & ~n_12176;
assign n_12178 =  x_1042 & ~n_12033;
assign n_12179 =  x_402 &  n_12033;
assign n_12180 = ~n_12178 & ~n_12179;
assign n_12181 =  x_1042 & ~n_12180;
assign n_12182 = ~x_1042 &  n_12180;
assign n_12183 = ~n_12181 & ~n_12182;
assign n_12184 =  x_1041 & ~n_12033;
assign n_12185 =  x_401 &  n_12033;
assign n_12186 = ~n_12184 & ~n_12185;
assign n_12187 =  x_1041 & ~n_12186;
assign n_12188 = ~x_1041 &  n_12186;
assign n_12189 = ~n_12187 & ~n_12188;
assign n_12190 =  x_1040 & ~n_12033;
assign n_12191 =  x_400 &  n_12033;
assign n_12192 = ~n_12190 & ~n_12191;
assign n_12193 =  x_1040 & ~n_12192;
assign n_12194 = ~x_1040 &  n_12192;
assign n_12195 = ~n_12193 & ~n_12194;
assign n_12196 =  x_1039 & ~n_12033;
assign n_12197 =  x_399 &  n_12033;
assign n_12198 = ~n_12196 & ~n_12197;
assign n_12199 =  x_1039 & ~n_12198;
assign n_12200 = ~x_1039 &  n_12198;
assign n_12201 = ~n_12199 & ~n_12200;
assign n_12202 =  x_1038 & ~n_12033;
assign n_12203 =  x_398 &  n_12033;
assign n_12204 = ~n_12202 & ~n_12203;
assign n_12205 =  x_1038 & ~n_12204;
assign n_12206 = ~x_1038 &  n_12204;
assign n_12207 = ~n_12205 & ~n_12206;
assign n_12208 =  x_1037 & ~n_12033;
assign n_12209 =  x_397 &  n_12033;
assign n_12210 = ~n_12208 & ~n_12209;
assign n_12211 =  x_1037 & ~n_12210;
assign n_12212 = ~x_1037 &  n_12210;
assign n_12213 = ~n_12211 & ~n_12212;
assign n_12214 =  x_1036 & ~n_12033;
assign n_12215 =  x_396 &  n_12033;
assign n_12216 = ~n_12214 & ~n_12215;
assign n_12217 =  x_1036 & ~n_12216;
assign n_12218 = ~x_1036 &  n_12216;
assign n_12219 = ~n_12217 & ~n_12218;
assign n_12220 =  x_1035 & ~n_12033;
assign n_12221 =  x_395 &  n_12033;
assign n_12222 = ~n_12220 & ~n_12221;
assign n_12223 =  x_1035 & ~n_12222;
assign n_12224 = ~x_1035 &  n_12222;
assign n_12225 = ~n_12223 & ~n_12224;
assign n_12226 = ~x_38 &  n_6330;
assign n_12227 =  n_3469 &  n_12226;
assign n_12228 =  x_1034 & ~n_12227;
assign n_12229 =  x_106 &  n_12227;
assign n_12230 = ~n_12228 & ~n_12229;
assign n_12231 =  x_1034 & ~n_12230;
assign n_12232 = ~x_1034 &  n_12230;
assign n_12233 = ~n_12231 & ~n_12232;
assign n_12234 =  x_1033 & ~n_12227;
assign n_12235 =  x_105 &  n_12227;
assign n_12236 = ~n_12234 & ~n_12235;
assign n_12237 =  x_1033 & ~n_12236;
assign n_12238 = ~x_1033 &  n_12236;
assign n_12239 = ~n_12237 & ~n_12238;
assign n_12240 =  x_1032 & ~n_12227;
assign n_12241 =  x_104 &  n_12227;
assign n_12242 = ~n_12240 & ~n_12241;
assign n_12243 =  x_1032 & ~n_12242;
assign n_12244 = ~x_1032 &  n_12242;
assign n_12245 = ~n_12243 & ~n_12244;
assign n_12246 =  x_1031 & ~n_12227;
assign n_12247 =  x_103 &  n_12227;
assign n_12248 = ~n_12246 & ~n_12247;
assign n_12249 =  x_1031 & ~n_12248;
assign n_12250 = ~x_1031 &  n_12248;
assign n_12251 = ~n_12249 & ~n_12250;
assign n_12252 =  x_1030 & ~n_12227;
assign n_12253 =  x_102 &  n_12227;
assign n_12254 = ~n_12252 & ~n_12253;
assign n_12255 =  x_1030 & ~n_12254;
assign n_12256 = ~x_1030 &  n_12254;
assign n_12257 = ~n_12255 & ~n_12256;
assign n_12258 =  x_1029 & ~n_12227;
assign n_12259 =  x_101 &  n_12227;
assign n_12260 = ~n_12258 & ~n_12259;
assign n_12261 =  x_1029 & ~n_12260;
assign n_12262 = ~x_1029 &  n_12260;
assign n_12263 = ~n_12261 & ~n_12262;
assign n_12264 =  x_1028 & ~n_12227;
assign n_12265 =  x_100 &  n_12227;
assign n_12266 = ~n_12264 & ~n_12265;
assign n_12267 =  x_1028 & ~n_12266;
assign n_12268 = ~x_1028 &  n_12266;
assign n_12269 = ~n_12267 & ~n_12268;
assign n_12270 =  x_1027 & ~n_12227;
assign n_12271 =  x_99 &  n_12227;
assign n_12272 = ~n_12270 & ~n_12271;
assign n_12273 =  x_1027 & ~n_12272;
assign n_12274 = ~x_1027 &  n_12272;
assign n_12275 = ~n_12273 & ~n_12274;
assign n_12276 =  x_1026 & ~n_12227;
assign n_12277 =  x_98 &  n_12227;
assign n_12278 = ~n_12276 & ~n_12277;
assign n_12279 =  x_1026 & ~n_12278;
assign n_12280 = ~x_1026 &  n_12278;
assign n_12281 = ~n_12279 & ~n_12280;
assign n_12282 =  x_1025 & ~n_12227;
assign n_12283 =  x_97 &  n_12227;
assign n_12284 = ~n_12282 & ~n_12283;
assign n_12285 =  x_1025 & ~n_12284;
assign n_12286 = ~x_1025 &  n_12284;
assign n_12287 = ~n_12285 & ~n_12286;
assign n_12288 =  x_1024 & ~n_12227;
assign n_12289 =  x_96 &  n_12227;
assign n_12290 = ~n_12288 & ~n_12289;
assign n_12291 =  x_1024 & ~n_12290;
assign n_12292 = ~x_1024 &  n_12290;
assign n_12293 = ~n_12291 & ~n_12292;
assign n_12294 =  x_1023 & ~n_12227;
assign n_12295 =  x_95 &  n_12227;
assign n_12296 = ~n_12294 & ~n_12295;
assign n_12297 =  x_1023 & ~n_12296;
assign n_12298 = ~x_1023 &  n_12296;
assign n_12299 = ~n_12297 & ~n_12298;
assign n_12300 =  x_1022 & ~n_12227;
assign n_12301 =  x_94 &  n_12227;
assign n_12302 = ~n_12300 & ~n_12301;
assign n_12303 =  x_1022 & ~n_12302;
assign n_12304 = ~x_1022 &  n_12302;
assign n_12305 = ~n_12303 & ~n_12304;
assign n_12306 =  x_1021 & ~n_12227;
assign n_12307 =  x_93 &  n_12227;
assign n_12308 = ~n_12306 & ~n_12307;
assign n_12309 =  x_1021 & ~n_12308;
assign n_12310 = ~x_1021 &  n_12308;
assign n_12311 = ~n_12309 & ~n_12310;
assign n_12312 =  x_1020 & ~n_12227;
assign n_12313 =  x_92 &  n_12227;
assign n_12314 = ~n_12312 & ~n_12313;
assign n_12315 =  x_1020 & ~n_12314;
assign n_12316 = ~x_1020 &  n_12314;
assign n_12317 = ~n_12315 & ~n_12316;
assign n_12318 =  x_1019 & ~n_12227;
assign n_12319 =  x_91 &  n_12227;
assign n_12320 = ~n_12318 & ~n_12319;
assign n_12321 =  x_1019 & ~n_12320;
assign n_12322 = ~x_1019 &  n_12320;
assign n_12323 = ~n_12321 & ~n_12322;
assign n_12324 =  x_1018 & ~n_12227;
assign n_12325 =  x_90 &  n_12227;
assign n_12326 = ~n_12324 & ~n_12325;
assign n_12327 =  x_1018 & ~n_12326;
assign n_12328 = ~x_1018 &  n_12326;
assign n_12329 = ~n_12327 & ~n_12328;
assign n_12330 =  x_1017 & ~n_12227;
assign n_12331 =  x_89 &  n_12227;
assign n_12332 = ~n_12330 & ~n_12331;
assign n_12333 =  x_1017 & ~n_12332;
assign n_12334 = ~x_1017 &  n_12332;
assign n_12335 = ~n_12333 & ~n_12334;
assign n_12336 =  x_1016 & ~n_12227;
assign n_12337 =  x_88 &  n_12227;
assign n_12338 = ~n_12336 & ~n_12337;
assign n_12339 =  x_1016 & ~n_12338;
assign n_12340 = ~x_1016 &  n_12338;
assign n_12341 = ~n_12339 & ~n_12340;
assign n_12342 =  x_1015 & ~n_12227;
assign n_12343 =  x_87 &  n_12227;
assign n_12344 = ~n_12342 & ~n_12343;
assign n_12345 =  x_1015 & ~n_12344;
assign n_12346 = ~x_1015 &  n_12344;
assign n_12347 = ~n_12345 & ~n_12346;
assign n_12348 =  x_1014 & ~n_12227;
assign n_12349 =  x_86 &  n_12227;
assign n_12350 = ~n_12348 & ~n_12349;
assign n_12351 =  x_1014 & ~n_12350;
assign n_12352 = ~x_1014 &  n_12350;
assign n_12353 = ~n_12351 & ~n_12352;
assign n_12354 =  x_1013 & ~n_12227;
assign n_12355 =  x_85 &  n_12227;
assign n_12356 = ~n_12354 & ~n_12355;
assign n_12357 =  x_1013 & ~n_12356;
assign n_12358 = ~x_1013 &  n_12356;
assign n_12359 = ~n_12357 & ~n_12358;
assign n_12360 =  x_1012 & ~n_12227;
assign n_12361 =  x_84 &  n_12227;
assign n_12362 = ~n_12360 & ~n_12361;
assign n_12363 =  x_1012 & ~n_12362;
assign n_12364 = ~x_1012 &  n_12362;
assign n_12365 = ~n_12363 & ~n_12364;
assign n_12366 =  x_1011 & ~n_12227;
assign n_12367 =  x_83 &  n_12227;
assign n_12368 = ~n_12366 & ~n_12367;
assign n_12369 =  x_1011 & ~n_12368;
assign n_12370 = ~x_1011 &  n_12368;
assign n_12371 = ~n_12369 & ~n_12370;
assign n_12372 =  x_1010 & ~n_12227;
assign n_12373 =  x_82 &  n_12227;
assign n_12374 = ~n_12372 & ~n_12373;
assign n_12375 =  x_1010 & ~n_12374;
assign n_12376 = ~x_1010 &  n_12374;
assign n_12377 = ~n_12375 & ~n_12376;
assign n_12378 =  x_1009 & ~n_12227;
assign n_12379 =  x_81 &  n_12227;
assign n_12380 = ~n_12378 & ~n_12379;
assign n_12381 =  x_1009 & ~n_12380;
assign n_12382 = ~x_1009 &  n_12380;
assign n_12383 = ~n_12381 & ~n_12382;
assign n_12384 =  x_1008 & ~n_12227;
assign n_12385 =  x_80 &  n_12227;
assign n_12386 = ~n_12384 & ~n_12385;
assign n_12387 =  x_1008 & ~n_12386;
assign n_12388 = ~x_1008 &  n_12386;
assign n_12389 = ~n_12387 & ~n_12388;
assign n_12390 =  x_1007 & ~n_12227;
assign n_12391 =  x_79 &  n_12227;
assign n_12392 = ~n_12390 & ~n_12391;
assign n_12393 =  x_1007 & ~n_12392;
assign n_12394 = ~x_1007 &  n_12392;
assign n_12395 = ~n_12393 & ~n_12394;
assign n_12396 =  x_1006 & ~n_12227;
assign n_12397 =  x_78 &  n_12227;
assign n_12398 = ~n_12396 & ~n_12397;
assign n_12399 =  x_1006 & ~n_12398;
assign n_12400 = ~x_1006 &  n_12398;
assign n_12401 = ~n_12399 & ~n_12400;
assign n_12402 =  x_1005 & ~n_12227;
assign n_12403 =  x_77 &  n_12227;
assign n_12404 = ~n_12402 & ~n_12403;
assign n_12405 =  x_1005 & ~n_12404;
assign n_12406 = ~x_1005 &  n_12404;
assign n_12407 = ~n_12405 & ~n_12406;
assign n_12408 =  x_1004 & ~n_12227;
assign n_12409 =  x_76 &  n_12227;
assign n_12410 = ~n_12408 & ~n_12409;
assign n_12411 =  x_1004 & ~n_12410;
assign n_12412 = ~x_1004 &  n_12410;
assign n_12413 = ~n_12411 & ~n_12412;
assign n_12414 =  x_1003 & ~n_12227;
assign n_12415 =  x_75 &  n_12227;
assign n_12416 = ~n_12414 & ~n_12415;
assign n_12417 =  x_1003 & ~n_12416;
assign n_12418 = ~x_1003 &  n_12416;
assign n_12419 = ~n_12417 & ~n_12418;
assign n_12420 =  n_4992 &  n_782;
assign n_12421 =  n_12420 &  n_4445;
assign n_12422 =  x_1002 & ~n_12421;
assign n_12423 =  i_32 &  n_12421;
assign n_12424 = ~n_12422 & ~n_12423;
assign n_12425 =  x_1002 & ~n_12424;
assign n_12426 = ~x_1002 &  n_12424;
assign n_12427 = ~n_12425 & ~n_12426;
assign n_12428 =  x_1001 & ~n_12421;
assign n_12429 =  i_31 &  n_12421;
assign n_12430 = ~n_12428 & ~n_12429;
assign n_12431 =  x_1001 & ~n_12430;
assign n_12432 = ~x_1001 &  n_12430;
assign n_12433 = ~n_12431 & ~n_12432;
assign n_12434 =  x_1000 & ~n_12421;
assign n_12435 =  i_30 &  n_12421;
assign n_12436 = ~n_12434 & ~n_12435;
assign n_12437 =  x_1000 & ~n_12436;
assign n_12438 = ~x_1000 &  n_12436;
assign n_12439 = ~n_12437 & ~n_12438;
assign n_12440 =  x_999 & ~n_12421;
assign n_12441 =  i_29 &  n_12421;
assign n_12442 = ~n_12440 & ~n_12441;
assign n_12443 =  x_999 & ~n_12442;
assign n_12444 = ~x_999 &  n_12442;
assign n_12445 = ~n_12443 & ~n_12444;
assign n_12446 =  x_998 & ~n_12421;
assign n_12447 =  i_28 &  n_12421;
assign n_12448 = ~n_12446 & ~n_12447;
assign n_12449 =  x_998 & ~n_12448;
assign n_12450 = ~x_998 &  n_12448;
assign n_12451 = ~n_12449 & ~n_12450;
assign n_12452 =  x_997 & ~n_12421;
assign n_12453 =  i_27 &  n_12421;
assign n_12454 = ~n_12452 & ~n_12453;
assign n_12455 =  x_997 & ~n_12454;
assign n_12456 = ~x_997 &  n_12454;
assign n_12457 = ~n_12455 & ~n_12456;
assign n_12458 =  x_996 & ~n_12421;
assign n_12459 =  i_26 &  n_12421;
assign n_12460 = ~n_12458 & ~n_12459;
assign n_12461 =  x_996 & ~n_12460;
assign n_12462 = ~x_996 &  n_12460;
assign n_12463 = ~n_12461 & ~n_12462;
assign n_12464 =  x_995 & ~n_12421;
assign n_12465 =  i_25 &  n_12421;
assign n_12466 = ~n_12464 & ~n_12465;
assign n_12467 =  x_995 & ~n_12466;
assign n_12468 = ~x_995 &  n_12466;
assign n_12469 = ~n_12467 & ~n_12468;
assign n_12470 =  x_994 & ~n_12421;
assign n_12471 =  i_24 &  n_12421;
assign n_12472 = ~n_12470 & ~n_12471;
assign n_12473 =  x_994 & ~n_12472;
assign n_12474 = ~x_994 &  n_12472;
assign n_12475 = ~n_12473 & ~n_12474;
assign n_12476 =  x_993 & ~n_12421;
assign n_12477 =  i_23 &  n_12421;
assign n_12478 = ~n_12476 & ~n_12477;
assign n_12479 =  x_993 & ~n_12478;
assign n_12480 = ~x_993 &  n_12478;
assign n_12481 = ~n_12479 & ~n_12480;
assign n_12482 =  x_992 & ~n_12421;
assign n_12483 =  i_22 &  n_12421;
assign n_12484 = ~n_12482 & ~n_12483;
assign n_12485 =  x_992 & ~n_12484;
assign n_12486 = ~x_992 &  n_12484;
assign n_12487 = ~n_12485 & ~n_12486;
assign n_12488 =  x_991 & ~n_12421;
assign n_12489 =  i_21 &  n_12421;
assign n_12490 = ~n_12488 & ~n_12489;
assign n_12491 =  x_991 & ~n_12490;
assign n_12492 = ~x_991 &  n_12490;
assign n_12493 = ~n_12491 & ~n_12492;
assign n_12494 =  x_990 & ~n_12421;
assign n_12495 =  i_20 &  n_12421;
assign n_12496 = ~n_12494 & ~n_12495;
assign n_12497 =  x_990 & ~n_12496;
assign n_12498 = ~x_990 &  n_12496;
assign n_12499 = ~n_12497 & ~n_12498;
assign n_12500 =  x_989 & ~n_12421;
assign n_12501 =  i_19 &  n_12421;
assign n_12502 = ~n_12500 & ~n_12501;
assign n_12503 =  x_989 & ~n_12502;
assign n_12504 = ~x_989 &  n_12502;
assign n_12505 = ~n_12503 & ~n_12504;
assign n_12506 =  x_988 & ~n_12421;
assign n_12507 =  i_18 &  n_12421;
assign n_12508 = ~n_12506 & ~n_12507;
assign n_12509 =  x_988 & ~n_12508;
assign n_12510 = ~x_988 &  n_12508;
assign n_12511 = ~n_12509 & ~n_12510;
assign n_12512 =  x_987 & ~n_12421;
assign n_12513 =  i_17 &  n_12421;
assign n_12514 = ~n_12512 & ~n_12513;
assign n_12515 =  x_987 & ~n_12514;
assign n_12516 = ~x_987 &  n_12514;
assign n_12517 = ~n_12515 & ~n_12516;
assign n_12518 =  x_986 & ~n_12421;
assign n_12519 =  i_16 &  n_12421;
assign n_12520 = ~n_12518 & ~n_12519;
assign n_12521 =  x_986 & ~n_12520;
assign n_12522 = ~x_986 &  n_12520;
assign n_12523 = ~n_12521 & ~n_12522;
assign n_12524 =  x_985 & ~n_12421;
assign n_12525 =  i_15 &  n_12421;
assign n_12526 = ~n_12524 & ~n_12525;
assign n_12527 =  x_985 & ~n_12526;
assign n_12528 = ~x_985 &  n_12526;
assign n_12529 = ~n_12527 & ~n_12528;
assign n_12530 =  x_984 & ~n_12421;
assign n_12531 =  i_14 &  n_12421;
assign n_12532 = ~n_12530 & ~n_12531;
assign n_12533 =  x_984 & ~n_12532;
assign n_12534 = ~x_984 &  n_12532;
assign n_12535 = ~n_12533 & ~n_12534;
assign n_12536 =  x_983 & ~n_12421;
assign n_12537 =  i_13 &  n_12421;
assign n_12538 = ~n_12536 & ~n_12537;
assign n_12539 =  x_983 & ~n_12538;
assign n_12540 = ~x_983 &  n_12538;
assign n_12541 = ~n_12539 & ~n_12540;
assign n_12542 =  x_982 & ~n_12421;
assign n_12543 =  i_12 &  n_12421;
assign n_12544 = ~n_12542 & ~n_12543;
assign n_12545 =  x_982 & ~n_12544;
assign n_12546 = ~x_982 &  n_12544;
assign n_12547 = ~n_12545 & ~n_12546;
assign n_12548 =  x_981 & ~n_12421;
assign n_12549 =  i_11 &  n_12421;
assign n_12550 = ~n_12548 & ~n_12549;
assign n_12551 =  x_981 & ~n_12550;
assign n_12552 = ~x_981 &  n_12550;
assign n_12553 = ~n_12551 & ~n_12552;
assign n_12554 =  x_980 & ~n_12421;
assign n_12555 =  i_10 &  n_12421;
assign n_12556 = ~n_12554 & ~n_12555;
assign n_12557 =  x_980 & ~n_12556;
assign n_12558 = ~x_980 &  n_12556;
assign n_12559 = ~n_12557 & ~n_12558;
assign n_12560 =  x_979 & ~n_12421;
assign n_12561 =  i_9 &  n_12421;
assign n_12562 = ~n_12560 & ~n_12561;
assign n_12563 =  x_979 & ~n_12562;
assign n_12564 = ~x_979 &  n_12562;
assign n_12565 = ~n_12563 & ~n_12564;
assign n_12566 =  x_978 & ~n_12421;
assign n_12567 =  i_8 &  n_12421;
assign n_12568 = ~n_12566 & ~n_12567;
assign n_12569 =  x_978 & ~n_12568;
assign n_12570 = ~x_978 &  n_12568;
assign n_12571 = ~n_12569 & ~n_12570;
assign n_12572 =  x_977 & ~n_12421;
assign n_12573 =  i_7 &  n_12421;
assign n_12574 = ~n_12572 & ~n_12573;
assign n_12575 =  x_977 & ~n_12574;
assign n_12576 = ~x_977 &  n_12574;
assign n_12577 = ~n_12575 & ~n_12576;
assign n_12578 =  x_976 & ~n_12421;
assign n_12579 =  i_6 &  n_12421;
assign n_12580 = ~n_12578 & ~n_12579;
assign n_12581 =  x_976 & ~n_12580;
assign n_12582 = ~x_976 &  n_12580;
assign n_12583 = ~n_12581 & ~n_12582;
assign n_12584 =  x_975 & ~n_12421;
assign n_12585 =  i_5 &  n_12421;
assign n_12586 = ~n_12584 & ~n_12585;
assign n_12587 =  x_975 & ~n_12586;
assign n_12588 = ~x_975 &  n_12586;
assign n_12589 = ~n_12587 & ~n_12588;
assign n_12590 =  x_974 & ~n_12421;
assign n_12591 =  i_4 &  n_12421;
assign n_12592 = ~n_12590 & ~n_12591;
assign n_12593 =  x_974 & ~n_12592;
assign n_12594 = ~x_974 &  n_12592;
assign n_12595 = ~n_12593 & ~n_12594;
assign n_12596 =  x_973 & ~n_12421;
assign n_12597 =  i_3 &  n_12421;
assign n_12598 = ~n_12596 & ~n_12597;
assign n_12599 =  x_973 & ~n_12598;
assign n_12600 = ~x_973 &  n_12598;
assign n_12601 = ~n_12599 & ~n_12600;
assign n_12602 =  x_972 & ~n_12421;
assign n_12603 =  i_2 &  n_12421;
assign n_12604 = ~n_12602 & ~n_12603;
assign n_12605 =  x_972 & ~n_12604;
assign n_12606 = ~x_972 &  n_12604;
assign n_12607 = ~n_12605 & ~n_12606;
assign n_12608 =  x_971 & ~n_12421;
assign n_12609 =  i_1 &  n_12421;
assign n_12610 = ~n_12608 & ~n_12609;
assign n_12611 =  x_971 & ~n_12610;
assign n_12612 = ~x_971 &  n_12610;
assign n_12613 = ~n_12611 & ~n_12612;
assign n_12614 = ~x_42 &  n_585;
assign n_12615 = ~x_39 &  n_4445;
assign n_12616 =  n_12614 &  n_12615;
assign n_12617 =  x_970 & ~n_12616;
assign n_12618 =  i_32 &  n_12616;
assign n_12619 = ~n_12617 & ~n_12618;
assign n_12620 =  x_970 & ~n_12619;
assign n_12621 = ~x_970 &  n_12619;
assign n_12622 = ~n_12620 & ~n_12621;
assign n_12623 =  x_969 & ~n_12616;
assign n_12624 =  i_31 &  n_12616;
assign n_12625 = ~n_12623 & ~n_12624;
assign n_12626 =  x_969 & ~n_12625;
assign n_12627 = ~x_969 &  n_12625;
assign n_12628 = ~n_12626 & ~n_12627;
assign n_12629 =  x_968 & ~n_12616;
assign n_12630 =  i_30 &  n_12616;
assign n_12631 = ~n_12629 & ~n_12630;
assign n_12632 =  x_968 & ~n_12631;
assign n_12633 = ~x_968 &  n_12631;
assign n_12634 = ~n_12632 & ~n_12633;
assign n_12635 =  x_967 & ~n_12616;
assign n_12636 =  i_29 &  n_12616;
assign n_12637 = ~n_12635 & ~n_12636;
assign n_12638 =  x_967 & ~n_12637;
assign n_12639 = ~x_967 &  n_12637;
assign n_12640 = ~n_12638 & ~n_12639;
assign n_12641 =  x_966 & ~n_12616;
assign n_12642 =  i_28 &  n_12616;
assign n_12643 = ~n_12641 & ~n_12642;
assign n_12644 =  x_966 & ~n_12643;
assign n_12645 = ~x_966 &  n_12643;
assign n_12646 = ~n_12644 & ~n_12645;
assign n_12647 =  x_965 & ~n_12616;
assign n_12648 =  i_27 &  n_12616;
assign n_12649 = ~n_12647 & ~n_12648;
assign n_12650 =  x_965 & ~n_12649;
assign n_12651 = ~x_965 &  n_12649;
assign n_12652 = ~n_12650 & ~n_12651;
assign n_12653 =  x_964 & ~n_12616;
assign n_12654 =  i_26 &  n_12616;
assign n_12655 = ~n_12653 & ~n_12654;
assign n_12656 =  x_964 & ~n_12655;
assign n_12657 = ~x_964 &  n_12655;
assign n_12658 = ~n_12656 & ~n_12657;
assign n_12659 =  x_963 & ~n_12616;
assign n_12660 =  i_25 &  n_12616;
assign n_12661 = ~n_12659 & ~n_12660;
assign n_12662 =  x_963 & ~n_12661;
assign n_12663 = ~x_963 &  n_12661;
assign n_12664 = ~n_12662 & ~n_12663;
assign n_12665 =  x_962 & ~n_12616;
assign n_12666 =  i_24 &  n_12616;
assign n_12667 = ~n_12665 & ~n_12666;
assign n_12668 =  x_962 & ~n_12667;
assign n_12669 = ~x_962 &  n_12667;
assign n_12670 = ~n_12668 & ~n_12669;
assign n_12671 =  x_961 & ~n_12616;
assign n_12672 =  i_23 &  n_12616;
assign n_12673 = ~n_12671 & ~n_12672;
assign n_12674 =  x_961 & ~n_12673;
assign n_12675 = ~x_961 &  n_12673;
assign n_12676 = ~n_12674 & ~n_12675;
assign n_12677 =  x_960 & ~n_12616;
assign n_12678 =  i_22 &  n_12616;
assign n_12679 = ~n_12677 & ~n_12678;
assign n_12680 =  x_960 & ~n_12679;
assign n_12681 = ~x_960 &  n_12679;
assign n_12682 = ~n_12680 & ~n_12681;
assign n_12683 =  x_959 & ~n_12616;
assign n_12684 =  i_21 &  n_12616;
assign n_12685 = ~n_12683 & ~n_12684;
assign n_12686 =  x_959 & ~n_12685;
assign n_12687 = ~x_959 &  n_12685;
assign n_12688 = ~n_12686 & ~n_12687;
assign n_12689 =  x_958 & ~n_12616;
assign n_12690 =  i_20 &  n_12616;
assign n_12691 = ~n_12689 & ~n_12690;
assign n_12692 =  x_958 & ~n_12691;
assign n_12693 = ~x_958 &  n_12691;
assign n_12694 = ~n_12692 & ~n_12693;
assign n_12695 =  x_957 & ~n_12616;
assign n_12696 =  i_19 &  n_12616;
assign n_12697 = ~n_12695 & ~n_12696;
assign n_12698 =  x_957 & ~n_12697;
assign n_12699 = ~x_957 &  n_12697;
assign n_12700 = ~n_12698 & ~n_12699;
assign n_12701 =  x_956 & ~n_12616;
assign n_12702 =  i_18 &  n_12616;
assign n_12703 = ~n_12701 & ~n_12702;
assign n_12704 =  x_956 & ~n_12703;
assign n_12705 = ~x_956 &  n_12703;
assign n_12706 = ~n_12704 & ~n_12705;
assign n_12707 =  x_955 & ~n_12616;
assign n_12708 =  i_17 &  n_12616;
assign n_12709 = ~n_12707 & ~n_12708;
assign n_12710 =  x_955 & ~n_12709;
assign n_12711 = ~x_955 &  n_12709;
assign n_12712 = ~n_12710 & ~n_12711;
assign n_12713 =  x_954 & ~n_12616;
assign n_12714 =  i_16 &  n_12616;
assign n_12715 = ~n_12713 & ~n_12714;
assign n_12716 =  x_954 & ~n_12715;
assign n_12717 = ~x_954 &  n_12715;
assign n_12718 = ~n_12716 & ~n_12717;
assign n_12719 =  x_953 & ~n_12616;
assign n_12720 =  i_15 &  n_12616;
assign n_12721 = ~n_12719 & ~n_12720;
assign n_12722 =  x_953 & ~n_12721;
assign n_12723 = ~x_953 &  n_12721;
assign n_12724 = ~n_12722 & ~n_12723;
assign n_12725 =  x_952 & ~n_12616;
assign n_12726 =  i_14 &  n_12616;
assign n_12727 = ~n_12725 & ~n_12726;
assign n_12728 =  x_952 & ~n_12727;
assign n_12729 = ~x_952 &  n_12727;
assign n_12730 = ~n_12728 & ~n_12729;
assign n_12731 =  x_951 & ~n_12616;
assign n_12732 =  i_13 &  n_12616;
assign n_12733 = ~n_12731 & ~n_12732;
assign n_12734 =  x_951 & ~n_12733;
assign n_12735 = ~x_951 &  n_12733;
assign n_12736 = ~n_12734 & ~n_12735;
assign n_12737 =  x_950 & ~n_12616;
assign n_12738 =  i_12 &  n_12616;
assign n_12739 = ~n_12737 & ~n_12738;
assign n_12740 =  x_950 & ~n_12739;
assign n_12741 = ~x_950 &  n_12739;
assign n_12742 = ~n_12740 & ~n_12741;
assign n_12743 =  x_949 & ~n_12616;
assign n_12744 =  i_11 &  n_12616;
assign n_12745 = ~n_12743 & ~n_12744;
assign n_12746 =  x_949 & ~n_12745;
assign n_12747 = ~x_949 &  n_12745;
assign n_12748 = ~n_12746 & ~n_12747;
assign n_12749 =  x_948 & ~n_12616;
assign n_12750 =  i_10 &  n_12616;
assign n_12751 = ~n_12749 & ~n_12750;
assign n_12752 =  x_948 & ~n_12751;
assign n_12753 = ~x_948 &  n_12751;
assign n_12754 = ~n_12752 & ~n_12753;
assign n_12755 =  x_947 & ~n_12616;
assign n_12756 =  i_9 &  n_12616;
assign n_12757 = ~n_12755 & ~n_12756;
assign n_12758 =  x_947 & ~n_12757;
assign n_12759 = ~x_947 &  n_12757;
assign n_12760 = ~n_12758 & ~n_12759;
assign n_12761 =  x_946 & ~n_12616;
assign n_12762 =  i_8 &  n_12616;
assign n_12763 = ~n_12761 & ~n_12762;
assign n_12764 =  x_946 & ~n_12763;
assign n_12765 = ~x_946 &  n_12763;
assign n_12766 = ~n_12764 & ~n_12765;
assign n_12767 =  x_945 & ~n_12616;
assign n_12768 =  i_7 &  n_12616;
assign n_12769 = ~n_12767 & ~n_12768;
assign n_12770 =  x_945 & ~n_12769;
assign n_12771 = ~x_945 &  n_12769;
assign n_12772 = ~n_12770 & ~n_12771;
assign n_12773 =  x_944 & ~n_12616;
assign n_12774 =  i_6 &  n_12616;
assign n_12775 = ~n_12773 & ~n_12774;
assign n_12776 =  x_944 & ~n_12775;
assign n_12777 = ~x_944 &  n_12775;
assign n_12778 = ~n_12776 & ~n_12777;
assign n_12779 =  x_943 & ~n_12616;
assign n_12780 =  i_5 &  n_12616;
assign n_12781 = ~n_12779 & ~n_12780;
assign n_12782 =  x_943 & ~n_12781;
assign n_12783 = ~x_943 &  n_12781;
assign n_12784 = ~n_12782 & ~n_12783;
assign n_12785 =  x_942 & ~n_12616;
assign n_12786 =  i_4 &  n_12616;
assign n_12787 = ~n_12785 & ~n_12786;
assign n_12788 =  x_942 & ~n_12787;
assign n_12789 = ~x_942 &  n_12787;
assign n_12790 = ~n_12788 & ~n_12789;
assign n_12791 =  x_941 & ~n_12616;
assign n_12792 =  i_3 &  n_12616;
assign n_12793 = ~n_12791 & ~n_12792;
assign n_12794 =  x_941 & ~n_12793;
assign n_12795 = ~x_941 &  n_12793;
assign n_12796 = ~n_12794 & ~n_12795;
assign n_12797 =  x_940 & ~n_12616;
assign n_12798 =  i_2 &  n_12616;
assign n_12799 = ~n_12797 & ~n_12798;
assign n_12800 =  x_940 & ~n_12799;
assign n_12801 = ~x_940 &  n_12799;
assign n_12802 = ~n_12800 & ~n_12801;
assign n_12803 =  x_939 & ~n_12616;
assign n_12804 =  i_1 &  n_12616;
assign n_12805 = ~n_12803 & ~n_12804;
assign n_12806 =  x_939 & ~n_12805;
assign n_12807 = ~x_939 &  n_12805;
assign n_12808 = ~n_12806 & ~n_12807;
assign n_12809 =  n_2 &  n_12615;
assign n_12810 =  x_938 & ~n_12809;
assign n_12811 =  i_32 &  n_12809;
assign n_12812 = ~n_12810 & ~n_12811;
assign n_12813 =  x_938 & ~n_12812;
assign n_12814 = ~x_938 &  n_12812;
assign n_12815 = ~n_12813 & ~n_12814;
assign n_12816 =  x_937 & ~n_12809;
assign n_12817 =  i_31 &  n_12809;
assign n_12818 = ~n_12816 & ~n_12817;
assign n_12819 =  x_937 & ~n_12818;
assign n_12820 = ~x_937 &  n_12818;
assign n_12821 = ~n_12819 & ~n_12820;
assign n_12822 =  x_936 & ~n_12809;
assign n_12823 =  i_30 &  n_12809;
assign n_12824 = ~n_12822 & ~n_12823;
assign n_12825 =  x_936 & ~n_12824;
assign n_12826 = ~x_936 &  n_12824;
assign n_12827 = ~n_12825 & ~n_12826;
assign n_12828 =  x_935 & ~n_12809;
assign n_12829 =  i_29 &  n_12809;
assign n_12830 = ~n_12828 & ~n_12829;
assign n_12831 =  x_935 & ~n_12830;
assign n_12832 = ~x_935 &  n_12830;
assign n_12833 = ~n_12831 & ~n_12832;
assign n_12834 =  x_934 & ~n_12809;
assign n_12835 =  i_28 &  n_12809;
assign n_12836 = ~n_12834 & ~n_12835;
assign n_12837 =  x_934 & ~n_12836;
assign n_12838 = ~x_934 &  n_12836;
assign n_12839 = ~n_12837 & ~n_12838;
assign n_12840 =  x_933 & ~n_12809;
assign n_12841 =  i_27 &  n_12809;
assign n_12842 = ~n_12840 & ~n_12841;
assign n_12843 =  x_933 & ~n_12842;
assign n_12844 = ~x_933 &  n_12842;
assign n_12845 = ~n_12843 & ~n_12844;
assign n_12846 =  x_932 & ~n_12809;
assign n_12847 =  i_26 &  n_12809;
assign n_12848 = ~n_12846 & ~n_12847;
assign n_12849 =  x_932 & ~n_12848;
assign n_12850 = ~x_932 &  n_12848;
assign n_12851 = ~n_12849 & ~n_12850;
assign n_12852 =  x_931 & ~n_12809;
assign n_12853 =  i_25 &  n_12809;
assign n_12854 = ~n_12852 & ~n_12853;
assign n_12855 =  x_931 & ~n_12854;
assign n_12856 = ~x_931 &  n_12854;
assign n_12857 = ~n_12855 & ~n_12856;
assign n_12858 =  x_930 & ~n_12809;
assign n_12859 =  i_24 &  n_12809;
assign n_12860 = ~n_12858 & ~n_12859;
assign n_12861 =  x_930 & ~n_12860;
assign n_12862 = ~x_930 &  n_12860;
assign n_12863 = ~n_12861 & ~n_12862;
assign n_12864 =  x_929 & ~n_12809;
assign n_12865 =  i_23 &  n_12809;
assign n_12866 = ~n_12864 & ~n_12865;
assign n_12867 =  x_929 & ~n_12866;
assign n_12868 = ~x_929 &  n_12866;
assign n_12869 = ~n_12867 & ~n_12868;
assign n_12870 =  x_928 & ~n_12809;
assign n_12871 =  i_22 &  n_12809;
assign n_12872 = ~n_12870 & ~n_12871;
assign n_12873 =  x_928 & ~n_12872;
assign n_12874 = ~x_928 &  n_12872;
assign n_12875 = ~n_12873 & ~n_12874;
assign n_12876 =  x_927 & ~n_12809;
assign n_12877 =  i_21 &  n_12809;
assign n_12878 = ~n_12876 & ~n_12877;
assign n_12879 =  x_927 & ~n_12878;
assign n_12880 = ~x_927 &  n_12878;
assign n_12881 = ~n_12879 & ~n_12880;
assign n_12882 =  x_926 & ~n_12809;
assign n_12883 =  i_20 &  n_12809;
assign n_12884 = ~n_12882 & ~n_12883;
assign n_12885 =  x_926 & ~n_12884;
assign n_12886 = ~x_926 &  n_12884;
assign n_12887 = ~n_12885 & ~n_12886;
assign n_12888 =  x_925 & ~n_12809;
assign n_12889 =  i_19 &  n_12809;
assign n_12890 = ~n_12888 & ~n_12889;
assign n_12891 =  x_925 & ~n_12890;
assign n_12892 = ~x_925 &  n_12890;
assign n_12893 = ~n_12891 & ~n_12892;
assign n_12894 =  x_924 & ~n_12809;
assign n_12895 =  i_18 &  n_12809;
assign n_12896 = ~n_12894 & ~n_12895;
assign n_12897 =  x_924 & ~n_12896;
assign n_12898 = ~x_924 &  n_12896;
assign n_12899 = ~n_12897 & ~n_12898;
assign n_12900 =  x_923 & ~n_12809;
assign n_12901 =  i_17 &  n_12809;
assign n_12902 = ~n_12900 & ~n_12901;
assign n_12903 =  x_923 & ~n_12902;
assign n_12904 = ~x_923 &  n_12902;
assign n_12905 = ~n_12903 & ~n_12904;
assign n_12906 =  x_922 & ~n_12809;
assign n_12907 =  i_16 &  n_12809;
assign n_12908 = ~n_12906 & ~n_12907;
assign n_12909 =  x_922 & ~n_12908;
assign n_12910 = ~x_922 &  n_12908;
assign n_12911 = ~n_12909 & ~n_12910;
assign n_12912 =  x_921 & ~n_12809;
assign n_12913 =  i_15 &  n_12809;
assign n_12914 = ~n_12912 & ~n_12913;
assign n_12915 =  x_921 & ~n_12914;
assign n_12916 = ~x_921 &  n_12914;
assign n_12917 = ~n_12915 & ~n_12916;
assign n_12918 =  x_920 & ~n_12809;
assign n_12919 =  i_14 &  n_12809;
assign n_12920 = ~n_12918 & ~n_12919;
assign n_12921 =  x_920 & ~n_12920;
assign n_12922 = ~x_920 &  n_12920;
assign n_12923 = ~n_12921 & ~n_12922;
assign n_12924 =  x_919 & ~n_12809;
assign n_12925 =  i_13 &  n_12809;
assign n_12926 = ~n_12924 & ~n_12925;
assign n_12927 =  x_919 & ~n_12926;
assign n_12928 = ~x_919 &  n_12926;
assign n_12929 = ~n_12927 & ~n_12928;
assign n_12930 =  x_918 & ~n_12809;
assign n_12931 =  i_12 &  n_12809;
assign n_12932 = ~n_12930 & ~n_12931;
assign n_12933 =  x_918 & ~n_12932;
assign n_12934 = ~x_918 &  n_12932;
assign n_12935 = ~n_12933 & ~n_12934;
assign n_12936 =  x_917 & ~n_12809;
assign n_12937 =  i_11 &  n_12809;
assign n_12938 = ~n_12936 & ~n_12937;
assign n_12939 =  x_917 & ~n_12938;
assign n_12940 = ~x_917 &  n_12938;
assign n_12941 = ~n_12939 & ~n_12940;
assign n_12942 =  x_916 & ~n_12809;
assign n_12943 =  i_10 &  n_12809;
assign n_12944 = ~n_12942 & ~n_12943;
assign n_12945 =  x_916 & ~n_12944;
assign n_12946 = ~x_916 &  n_12944;
assign n_12947 = ~n_12945 & ~n_12946;
assign n_12948 =  x_915 & ~n_12809;
assign n_12949 =  i_9 &  n_12809;
assign n_12950 = ~n_12948 & ~n_12949;
assign n_12951 =  x_915 & ~n_12950;
assign n_12952 = ~x_915 &  n_12950;
assign n_12953 = ~n_12951 & ~n_12952;
assign n_12954 =  x_914 & ~n_12809;
assign n_12955 =  i_8 &  n_12809;
assign n_12956 = ~n_12954 & ~n_12955;
assign n_12957 =  x_914 & ~n_12956;
assign n_12958 = ~x_914 &  n_12956;
assign n_12959 = ~n_12957 & ~n_12958;
assign n_12960 =  x_913 & ~n_12809;
assign n_12961 =  i_7 &  n_12809;
assign n_12962 = ~n_12960 & ~n_12961;
assign n_12963 =  x_913 & ~n_12962;
assign n_12964 = ~x_913 &  n_12962;
assign n_12965 = ~n_12963 & ~n_12964;
assign n_12966 =  x_912 & ~n_12809;
assign n_12967 =  i_6 &  n_12809;
assign n_12968 = ~n_12966 & ~n_12967;
assign n_12969 =  x_912 & ~n_12968;
assign n_12970 = ~x_912 &  n_12968;
assign n_12971 = ~n_12969 & ~n_12970;
assign n_12972 =  x_911 & ~n_12809;
assign n_12973 =  i_5 &  n_12809;
assign n_12974 = ~n_12972 & ~n_12973;
assign n_12975 =  x_911 & ~n_12974;
assign n_12976 = ~x_911 &  n_12974;
assign n_12977 = ~n_12975 & ~n_12976;
assign n_12978 =  x_910 & ~n_12809;
assign n_12979 =  i_4 &  n_12809;
assign n_12980 = ~n_12978 & ~n_12979;
assign n_12981 =  x_910 & ~n_12980;
assign n_12982 = ~x_910 &  n_12980;
assign n_12983 = ~n_12981 & ~n_12982;
assign n_12984 =  x_909 & ~n_12809;
assign n_12985 =  i_3 &  n_12809;
assign n_12986 = ~n_12984 & ~n_12985;
assign n_12987 =  x_909 & ~n_12986;
assign n_12988 = ~x_909 &  n_12986;
assign n_12989 = ~n_12987 & ~n_12988;
assign n_12990 =  x_908 & ~n_12809;
assign n_12991 =  i_2 &  n_12809;
assign n_12992 = ~n_12990 & ~n_12991;
assign n_12993 =  x_908 & ~n_12992;
assign n_12994 = ~x_908 &  n_12992;
assign n_12995 = ~n_12993 & ~n_12994;
assign n_12996 =  x_907 & ~n_12809;
assign n_12997 =  i_1 &  n_12809;
assign n_12998 = ~n_12996 & ~n_12997;
assign n_12999 =  x_907 & ~n_12998;
assign n_13000 = ~x_907 &  n_12998;
assign n_13001 = ~n_12999 & ~n_13000;
assign n_13002 =  x_41 &  n_184;
assign n_13003 = ~n_4057 & ~n_7865;
assign n_13004 =  n_13002 & ~n_13003;
assign n_13005 =  x_39 &  n_1312;
assign n_13006 =  n_981 &  n_13005;
assign n_13007 = ~n_2301 &  n_13006;
assign n_13008 =  n_585 &  n_8803;
assign n_13009 = ~n_13007 & ~n_13008;
assign n_13010 = ~n_13004 &  n_13009;
assign n_13011 = ~x_42 & ~n_13010;
assign n_13012 =  x_42 &  n_2301;
assign n_13013 =  n_13012 &  n_4251;
assign n_13014 = ~x_42 &  n_2301;
assign n_13015 =  n_1313 &  n_981;
assign n_13016 =  n_13014 &  n_13015;
assign n_13017 = ~n_13013 & ~n_13016;
assign n_13018 = ~n_13011 &  n_13017;
assign n_13019 =  x_906 &  n_13018;
assign n_13020 =  n_184 &  n_7865;
assign n_13021 =  n_185 &  n_13020;
assign n_13022 = ~x_42 &  n_13007;
assign n_13023 = ~n_13021 & ~n_13022;
assign n_13024 =  i_32 & ~n_13023;
assign n_13025 =  n_185 &  n_10521;
assign n_13026 =  x_1098 &  n_13025;
assign n_13027 =  x_554 &  n_13013;
assign n_13028 = ~n_13026 & ~n_13027;
assign n_13029 =  x_522 &  n_13016;
assign n_13030 =  n_12614 &  n_8803;
assign n_13031 =  x_1162 &  n_13030;
assign n_13032 = ~n_13029 & ~n_13031;
assign n_13033 =  n_13028 &  n_13032;
assign n_13034 = ~n_13024 &  n_13033;
assign n_13035 = ~n_13019 &  n_13034;
assign n_13036 =  x_906 & ~n_13035;
assign n_13037 = ~x_906 &  n_13035;
assign n_13038 = ~n_13036 & ~n_13037;
assign n_13039 =  x_905 &  n_13018;
assign n_13040 =  i_31 & ~n_13023;
assign n_13041 =  x_1097 &  n_13025;
assign n_13042 =  x_553 &  n_13013;
assign n_13043 = ~n_13041 & ~n_13042;
assign n_13044 =  x_521 &  n_13016;
assign n_13045 =  x_1161 &  n_13030;
assign n_13046 = ~n_13044 & ~n_13045;
assign n_13047 =  n_13043 &  n_13046;
assign n_13048 = ~n_13040 &  n_13047;
assign n_13049 = ~n_13039 &  n_13048;
assign n_13050 =  x_905 & ~n_13049;
assign n_13051 = ~x_905 &  n_13049;
assign n_13052 = ~n_13050 & ~n_13051;
assign n_13053 =  x_904 &  n_13018;
assign n_13054 =  i_30 & ~n_13023;
assign n_13055 =  x_1096 &  n_13025;
assign n_13056 =  x_552 &  n_13013;
assign n_13057 = ~n_13055 & ~n_13056;
assign n_13058 =  x_520 &  n_13016;
assign n_13059 =  x_1160 &  n_13030;
assign n_13060 = ~n_13058 & ~n_13059;
assign n_13061 =  n_13057 &  n_13060;
assign n_13062 = ~n_13054 &  n_13061;
assign n_13063 = ~n_13053 &  n_13062;
assign n_13064 =  x_904 & ~n_13063;
assign n_13065 = ~x_904 &  n_13063;
assign n_13066 = ~n_13064 & ~n_13065;
assign n_13067 =  x_903 &  n_13018;
assign n_13068 =  i_29 & ~n_13023;
assign n_13069 =  x_1095 &  n_13025;
assign n_13070 =  x_551 &  n_13013;
assign n_13071 = ~n_13069 & ~n_13070;
assign n_13072 =  x_519 &  n_13016;
assign n_13073 =  x_1159 &  n_13030;
assign n_13074 = ~n_13072 & ~n_13073;
assign n_13075 =  n_13071 &  n_13074;
assign n_13076 = ~n_13068 &  n_13075;
assign n_13077 = ~n_13067 &  n_13076;
assign n_13078 =  x_903 & ~n_13077;
assign n_13079 = ~x_903 &  n_13077;
assign n_13080 = ~n_13078 & ~n_13079;
assign n_13081 =  x_902 &  n_13018;
assign n_13082 =  i_28 & ~n_13023;
assign n_13083 =  x_1094 &  n_13025;
assign n_13084 =  x_550 &  n_13013;
assign n_13085 = ~n_13083 & ~n_13084;
assign n_13086 =  x_518 &  n_13016;
assign n_13087 =  x_1158 &  n_13030;
assign n_13088 = ~n_13086 & ~n_13087;
assign n_13089 =  n_13085 &  n_13088;
assign n_13090 = ~n_13082 &  n_13089;
assign n_13091 = ~n_13081 &  n_13090;
assign n_13092 =  x_902 & ~n_13091;
assign n_13093 = ~x_902 &  n_13091;
assign n_13094 = ~n_13092 & ~n_13093;
assign n_13095 =  x_901 &  n_13018;
assign n_13096 =  i_27 & ~n_13023;
assign n_13097 =  x_1093 &  n_13025;
assign n_13098 =  x_549 &  n_13013;
assign n_13099 = ~n_13097 & ~n_13098;
assign n_13100 =  x_517 &  n_13016;
assign n_13101 =  x_1157 &  n_13030;
assign n_13102 = ~n_13100 & ~n_13101;
assign n_13103 =  n_13099 &  n_13102;
assign n_13104 = ~n_13096 &  n_13103;
assign n_13105 = ~n_13095 &  n_13104;
assign n_13106 =  x_901 & ~n_13105;
assign n_13107 = ~x_901 &  n_13105;
assign n_13108 = ~n_13106 & ~n_13107;
assign n_13109 =  x_900 &  n_13018;
assign n_13110 =  i_26 & ~n_13023;
assign n_13111 =  x_1092 &  n_13025;
assign n_13112 =  x_548 &  n_13013;
assign n_13113 = ~n_13111 & ~n_13112;
assign n_13114 =  x_516 &  n_13016;
assign n_13115 =  x_1156 &  n_13030;
assign n_13116 = ~n_13114 & ~n_13115;
assign n_13117 =  n_13113 &  n_13116;
assign n_13118 = ~n_13110 &  n_13117;
assign n_13119 = ~n_13109 &  n_13118;
assign n_13120 =  x_900 & ~n_13119;
assign n_13121 = ~x_900 &  n_13119;
assign n_13122 = ~n_13120 & ~n_13121;
assign n_13123 =  x_899 &  n_13018;
assign n_13124 =  i_25 & ~n_13023;
assign n_13125 =  x_1091 &  n_13025;
assign n_13126 =  x_547 &  n_13013;
assign n_13127 = ~n_13125 & ~n_13126;
assign n_13128 =  x_515 &  n_13016;
assign n_13129 =  x_1155 &  n_13030;
assign n_13130 = ~n_13128 & ~n_13129;
assign n_13131 =  n_13127 &  n_13130;
assign n_13132 = ~n_13124 &  n_13131;
assign n_13133 = ~n_13123 &  n_13132;
assign n_13134 =  x_899 & ~n_13133;
assign n_13135 = ~x_899 &  n_13133;
assign n_13136 = ~n_13134 & ~n_13135;
assign n_13137 =  x_898 &  n_13018;
assign n_13138 =  i_24 & ~n_13023;
assign n_13139 =  x_1090 &  n_13025;
assign n_13140 =  x_546 &  n_13013;
assign n_13141 = ~n_13139 & ~n_13140;
assign n_13142 =  x_514 &  n_13016;
assign n_13143 =  x_1154 &  n_13030;
assign n_13144 = ~n_13142 & ~n_13143;
assign n_13145 =  n_13141 &  n_13144;
assign n_13146 = ~n_13138 &  n_13145;
assign n_13147 = ~n_13137 &  n_13146;
assign n_13148 =  x_898 & ~n_13147;
assign n_13149 = ~x_898 &  n_13147;
assign n_13150 = ~n_13148 & ~n_13149;
assign n_13151 =  x_897 &  n_13018;
assign n_13152 =  i_23 & ~n_13023;
assign n_13153 =  x_1089 &  n_13025;
assign n_13154 =  x_545 &  n_13013;
assign n_13155 = ~n_13153 & ~n_13154;
assign n_13156 =  x_513 &  n_13016;
assign n_13157 =  x_1153 &  n_13030;
assign n_13158 = ~n_13156 & ~n_13157;
assign n_13159 =  n_13155 &  n_13158;
assign n_13160 = ~n_13152 &  n_13159;
assign n_13161 = ~n_13151 &  n_13160;
assign n_13162 =  x_897 & ~n_13161;
assign n_13163 = ~x_897 &  n_13161;
assign n_13164 = ~n_13162 & ~n_13163;
assign n_13165 =  x_896 &  n_13018;
assign n_13166 =  i_22 & ~n_13023;
assign n_13167 =  x_1088 &  n_13025;
assign n_13168 =  x_544 &  n_13013;
assign n_13169 = ~n_13167 & ~n_13168;
assign n_13170 =  x_512 &  n_13016;
assign n_13171 =  x_1152 &  n_13030;
assign n_13172 = ~n_13170 & ~n_13171;
assign n_13173 =  n_13169 &  n_13172;
assign n_13174 = ~n_13166 &  n_13173;
assign n_13175 = ~n_13165 &  n_13174;
assign n_13176 =  x_896 & ~n_13175;
assign n_13177 = ~x_896 &  n_13175;
assign n_13178 = ~n_13176 & ~n_13177;
assign n_13179 =  x_895 &  n_13018;
assign n_13180 =  i_21 & ~n_13023;
assign n_13181 =  x_1087 &  n_13025;
assign n_13182 =  x_543 &  n_13013;
assign n_13183 = ~n_13181 & ~n_13182;
assign n_13184 =  x_511 &  n_13016;
assign n_13185 =  x_1151 &  n_13030;
assign n_13186 = ~n_13184 & ~n_13185;
assign n_13187 =  n_13183 &  n_13186;
assign n_13188 = ~n_13180 &  n_13187;
assign n_13189 = ~n_13179 &  n_13188;
assign n_13190 =  x_895 & ~n_13189;
assign n_13191 = ~x_895 &  n_13189;
assign n_13192 = ~n_13190 & ~n_13191;
assign n_13193 =  x_894 &  n_13018;
assign n_13194 =  i_20 & ~n_13023;
assign n_13195 =  x_1086 &  n_13025;
assign n_13196 =  x_542 &  n_13013;
assign n_13197 = ~n_13195 & ~n_13196;
assign n_13198 =  x_510 &  n_13016;
assign n_13199 =  x_1150 &  n_13030;
assign n_13200 = ~n_13198 & ~n_13199;
assign n_13201 =  n_13197 &  n_13200;
assign n_13202 = ~n_13194 &  n_13201;
assign n_13203 = ~n_13193 &  n_13202;
assign n_13204 =  x_894 & ~n_13203;
assign n_13205 = ~x_894 &  n_13203;
assign n_13206 = ~n_13204 & ~n_13205;
assign n_13207 =  x_893 &  n_13018;
assign n_13208 =  i_19 & ~n_13023;
assign n_13209 =  x_1085 &  n_13025;
assign n_13210 =  x_541 &  n_13013;
assign n_13211 = ~n_13209 & ~n_13210;
assign n_13212 =  x_509 &  n_13016;
assign n_13213 =  x_1149 &  n_13030;
assign n_13214 = ~n_13212 & ~n_13213;
assign n_13215 =  n_13211 &  n_13214;
assign n_13216 = ~n_13208 &  n_13215;
assign n_13217 = ~n_13207 &  n_13216;
assign n_13218 =  x_893 & ~n_13217;
assign n_13219 = ~x_893 &  n_13217;
assign n_13220 = ~n_13218 & ~n_13219;
assign n_13221 =  x_892 &  n_13018;
assign n_13222 =  i_18 & ~n_13023;
assign n_13223 =  x_1084 &  n_13025;
assign n_13224 =  x_540 &  n_13013;
assign n_13225 = ~n_13223 & ~n_13224;
assign n_13226 =  x_508 &  n_13016;
assign n_13227 =  x_1148 &  n_13030;
assign n_13228 = ~n_13226 & ~n_13227;
assign n_13229 =  n_13225 &  n_13228;
assign n_13230 = ~n_13222 &  n_13229;
assign n_13231 = ~n_13221 &  n_13230;
assign n_13232 =  x_892 & ~n_13231;
assign n_13233 = ~x_892 &  n_13231;
assign n_13234 = ~n_13232 & ~n_13233;
assign n_13235 =  x_891 &  n_13018;
assign n_13236 =  i_17 & ~n_13023;
assign n_13237 =  x_1083 &  n_13025;
assign n_13238 =  x_539 &  n_13013;
assign n_13239 = ~n_13237 & ~n_13238;
assign n_13240 =  x_507 &  n_13016;
assign n_13241 =  x_1147 &  n_13030;
assign n_13242 = ~n_13240 & ~n_13241;
assign n_13243 =  n_13239 &  n_13242;
assign n_13244 = ~n_13236 &  n_13243;
assign n_13245 = ~n_13235 &  n_13244;
assign n_13246 =  x_891 & ~n_13245;
assign n_13247 = ~x_891 &  n_13245;
assign n_13248 = ~n_13246 & ~n_13247;
assign n_13249 =  x_890 &  n_13018;
assign n_13250 =  i_16 & ~n_13023;
assign n_13251 =  x_1082 &  n_13025;
assign n_13252 =  x_538 &  n_13013;
assign n_13253 = ~n_13251 & ~n_13252;
assign n_13254 =  x_506 &  n_13016;
assign n_13255 =  x_1146 &  n_13030;
assign n_13256 = ~n_13254 & ~n_13255;
assign n_13257 =  n_13253 &  n_13256;
assign n_13258 = ~n_13250 &  n_13257;
assign n_13259 = ~n_13249 &  n_13258;
assign n_13260 =  x_890 & ~n_13259;
assign n_13261 = ~x_890 &  n_13259;
assign n_13262 = ~n_13260 & ~n_13261;
assign n_13263 =  x_889 &  n_13018;
assign n_13264 =  i_15 & ~n_13023;
assign n_13265 =  x_1081 &  n_13025;
assign n_13266 =  x_537 &  n_13013;
assign n_13267 = ~n_13265 & ~n_13266;
assign n_13268 =  x_505 &  n_13016;
assign n_13269 =  x_1145 &  n_13030;
assign n_13270 = ~n_13268 & ~n_13269;
assign n_13271 =  n_13267 &  n_13270;
assign n_13272 = ~n_13264 &  n_13271;
assign n_13273 = ~n_13263 &  n_13272;
assign n_13274 =  x_889 & ~n_13273;
assign n_13275 = ~x_889 &  n_13273;
assign n_13276 = ~n_13274 & ~n_13275;
assign n_13277 =  x_888 &  n_13018;
assign n_13278 =  i_14 & ~n_13023;
assign n_13279 =  x_1080 &  n_13025;
assign n_13280 =  x_536 &  n_13013;
assign n_13281 = ~n_13279 & ~n_13280;
assign n_13282 =  x_504 &  n_13016;
assign n_13283 =  x_1144 &  n_13030;
assign n_13284 = ~n_13282 & ~n_13283;
assign n_13285 =  n_13281 &  n_13284;
assign n_13286 = ~n_13278 &  n_13285;
assign n_13287 = ~n_13277 &  n_13286;
assign n_13288 =  x_888 & ~n_13287;
assign n_13289 = ~x_888 &  n_13287;
assign n_13290 = ~n_13288 & ~n_13289;
assign n_13291 =  x_887 &  n_13018;
assign n_13292 =  i_13 & ~n_13023;
assign n_13293 =  x_1079 &  n_13025;
assign n_13294 =  x_535 &  n_13013;
assign n_13295 = ~n_13293 & ~n_13294;
assign n_13296 =  x_503 &  n_13016;
assign n_13297 =  x_1143 &  n_13030;
assign n_13298 = ~n_13296 & ~n_13297;
assign n_13299 =  n_13295 &  n_13298;
assign n_13300 = ~n_13292 &  n_13299;
assign n_13301 = ~n_13291 &  n_13300;
assign n_13302 =  x_887 & ~n_13301;
assign n_13303 = ~x_887 &  n_13301;
assign n_13304 = ~n_13302 & ~n_13303;
assign n_13305 =  x_886 &  n_13018;
assign n_13306 =  i_12 & ~n_13023;
assign n_13307 =  x_1078 &  n_13025;
assign n_13308 =  x_534 &  n_13013;
assign n_13309 = ~n_13307 & ~n_13308;
assign n_13310 =  x_502 &  n_13016;
assign n_13311 =  x_1142 &  n_13030;
assign n_13312 = ~n_13310 & ~n_13311;
assign n_13313 =  n_13309 &  n_13312;
assign n_13314 = ~n_13306 &  n_13313;
assign n_13315 = ~n_13305 &  n_13314;
assign n_13316 =  x_886 & ~n_13315;
assign n_13317 = ~x_886 &  n_13315;
assign n_13318 = ~n_13316 & ~n_13317;
assign n_13319 =  x_885 &  n_13018;
assign n_13320 =  i_11 & ~n_13023;
assign n_13321 =  x_1077 &  n_13025;
assign n_13322 =  x_533 &  n_13013;
assign n_13323 = ~n_13321 & ~n_13322;
assign n_13324 =  x_501 &  n_13016;
assign n_13325 =  x_1141 &  n_13030;
assign n_13326 = ~n_13324 & ~n_13325;
assign n_13327 =  n_13323 &  n_13326;
assign n_13328 = ~n_13320 &  n_13327;
assign n_13329 = ~n_13319 &  n_13328;
assign n_13330 =  x_885 & ~n_13329;
assign n_13331 = ~x_885 &  n_13329;
assign n_13332 = ~n_13330 & ~n_13331;
assign n_13333 =  x_884 &  n_13018;
assign n_13334 =  i_10 & ~n_13023;
assign n_13335 =  x_1076 &  n_13025;
assign n_13336 =  x_532 &  n_13013;
assign n_13337 = ~n_13335 & ~n_13336;
assign n_13338 =  x_500 &  n_13016;
assign n_13339 =  x_1140 &  n_13030;
assign n_13340 = ~n_13338 & ~n_13339;
assign n_13341 =  n_13337 &  n_13340;
assign n_13342 = ~n_13334 &  n_13341;
assign n_13343 = ~n_13333 &  n_13342;
assign n_13344 =  x_884 & ~n_13343;
assign n_13345 = ~x_884 &  n_13343;
assign n_13346 = ~n_13344 & ~n_13345;
assign n_13347 =  x_883 &  n_13018;
assign n_13348 =  i_9 & ~n_13023;
assign n_13349 =  x_1075 &  n_13025;
assign n_13350 =  x_531 &  n_13013;
assign n_13351 = ~n_13349 & ~n_13350;
assign n_13352 =  x_499 &  n_13016;
assign n_13353 =  x_1139 &  n_13030;
assign n_13354 = ~n_13352 & ~n_13353;
assign n_13355 =  n_13351 &  n_13354;
assign n_13356 = ~n_13348 &  n_13355;
assign n_13357 = ~n_13347 &  n_13356;
assign n_13358 =  x_883 & ~n_13357;
assign n_13359 = ~x_883 &  n_13357;
assign n_13360 = ~n_13358 & ~n_13359;
assign n_13361 =  x_882 &  n_13018;
assign n_13362 =  i_8 & ~n_13023;
assign n_13363 =  x_1074 &  n_13025;
assign n_13364 =  x_530 &  n_13013;
assign n_13365 = ~n_13363 & ~n_13364;
assign n_13366 =  x_498 &  n_13016;
assign n_13367 =  x_1138 &  n_13030;
assign n_13368 = ~n_13366 & ~n_13367;
assign n_13369 =  n_13365 &  n_13368;
assign n_13370 = ~n_13362 &  n_13369;
assign n_13371 = ~n_13361 &  n_13370;
assign n_13372 =  x_882 & ~n_13371;
assign n_13373 = ~x_882 &  n_13371;
assign n_13374 = ~n_13372 & ~n_13373;
assign n_13375 =  x_881 &  n_13018;
assign n_13376 =  i_7 & ~n_13023;
assign n_13377 =  x_1073 &  n_13025;
assign n_13378 =  x_529 &  n_13013;
assign n_13379 = ~n_13377 & ~n_13378;
assign n_13380 =  x_497 &  n_13016;
assign n_13381 =  x_1137 &  n_13030;
assign n_13382 = ~n_13380 & ~n_13381;
assign n_13383 =  n_13379 &  n_13382;
assign n_13384 = ~n_13376 &  n_13383;
assign n_13385 = ~n_13375 &  n_13384;
assign n_13386 =  x_881 & ~n_13385;
assign n_13387 = ~x_881 &  n_13385;
assign n_13388 = ~n_13386 & ~n_13387;
assign n_13389 =  x_880 &  n_13018;
assign n_13390 =  i_6 & ~n_13023;
assign n_13391 =  x_1072 &  n_13025;
assign n_13392 =  x_528 &  n_13013;
assign n_13393 = ~n_13391 & ~n_13392;
assign n_13394 =  x_496 &  n_13016;
assign n_13395 =  x_1136 &  n_13030;
assign n_13396 = ~n_13394 & ~n_13395;
assign n_13397 =  n_13393 &  n_13396;
assign n_13398 = ~n_13390 &  n_13397;
assign n_13399 = ~n_13389 &  n_13398;
assign n_13400 =  x_880 & ~n_13399;
assign n_13401 = ~x_880 &  n_13399;
assign n_13402 = ~n_13400 & ~n_13401;
assign n_13403 =  x_879 &  n_13018;
assign n_13404 =  i_5 & ~n_13023;
assign n_13405 =  x_1071 &  n_13025;
assign n_13406 =  x_527 &  n_13013;
assign n_13407 = ~n_13405 & ~n_13406;
assign n_13408 =  x_495 &  n_13016;
assign n_13409 =  x_1135 &  n_13030;
assign n_13410 = ~n_13408 & ~n_13409;
assign n_13411 =  n_13407 &  n_13410;
assign n_13412 = ~n_13404 &  n_13411;
assign n_13413 = ~n_13403 &  n_13412;
assign n_13414 =  x_879 & ~n_13413;
assign n_13415 = ~x_879 &  n_13413;
assign n_13416 = ~n_13414 & ~n_13415;
assign n_13417 =  x_878 &  n_13018;
assign n_13418 =  i_4 & ~n_13023;
assign n_13419 =  x_1070 &  n_13025;
assign n_13420 =  x_526 &  n_13013;
assign n_13421 = ~n_13419 & ~n_13420;
assign n_13422 =  x_494 &  n_13016;
assign n_13423 =  x_1134 &  n_13030;
assign n_13424 = ~n_13422 & ~n_13423;
assign n_13425 =  n_13421 &  n_13424;
assign n_13426 = ~n_13418 &  n_13425;
assign n_13427 = ~n_13417 &  n_13426;
assign n_13428 =  x_878 & ~n_13427;
assign n_13429 = ~x_878 &  n_13427;
assign n_13430 = ~n_13428 & ~n_13429;
assign n_13431 =  x_877 &  n_13018;
assign n_13432 =  i_3 & ~n_13023;
assign n_13433 =  x_1069 &  n_13025;
assign n_13434 =  x_525 &  n_13013;
assign n_13435 = ~n_13433 & ~n_13434;
assign n_13436 =  x_493 &  n_13016;
assign n_13437 =  x_1133 &  n_13030;
assign n_13438 = ~n_13436 & ~n_13437;
assign n_13439 =  n_13435 &  n_13438;
assign n_13440 = ~n_13432 &  n_13439;
assign n_13441 = ~n_13431 &  n_13440;
assign n_13442 =  x_877 & ~n_13441;
assign n_13443 = ~x_877 &  n_13441;
assign n_13444 = ~n_13442 & ~n_13443;
assign n_13445 =  x_876 &  n_13018;
assign n_13446 =  i_2 & ~n_13023;
assign n_13447 =  x_1068 &  n_13025;
assign n_13448 =  x_524 &  n_13013;
assign n_13449 = ~n_13447 & ~n_13448;
assign n_13450 =  x_492 &  n_13016;
assign n_13451 =  x_1132 &  n_13030;
assign n_13452 = ~n_13450 & ~n_13451;
assign n_13453 =  n_13449 &  n_13452;
assign n_13454 = ~n_13446 &  n_13453;
assign n_13455 = ~n_13445 &  n_13454;
assign n_13456 =  x_876 & ~n_13455;
assign n_13457 = ~x_876 &  n_13455;
assign n_13458 = ~n_13456 & ~n_13457;
assign n_13459 =  x_875 &  n_13018;
assign n_13460 =  i_1 & ~n_13023;
assign n_13461 =  x_1067 &  n_13025;
assign n_13462 =  x_523 &  n_13013;
assign n_13463 = ~n_13461 & ~n_13462;
assign n_13464 =  x_491 &  n_13016;
assign n_13465 =  x_1131 &  n_13030;
assign n_13466 = ~n_13464 & ~n_13465;
assign n_13467 =  n_13463 &  n_13466;
assign n_13468 = ~n_13460 &  n_13467;
assign n_13469 = ~n_13459 &  n_13468;
assign n_13470 =  x_875 & ~n_13469;
assign n_13471 = ~x_875 &  n_13469;
assign n_13472 = ~n_13470 & ~n_13471;
assign n_13473 =  n_1 &  n_10515;
assign n_13474 = ~x_42 &  n_13473;
assign n_13475 =  x_874 & ~n_13474;
assign n_13476 =  x_106 &  n_13474;
assign n_13477 = ~n_13475 & ~n_13476;
assign n_13478 =  x_874 & ~n_13477;
assign n_13479 = ~x_874 &  n_13477;
assign n_13480 = ~n_13478 & ~n_13479;
assign n_13481 =  x_873 & ~n_13474;
assign n_13482 =  x_105 &  n_13474;
assign n_13483 = ~n_13481 & ~n_13482;
assign n_13484 =  x_873 & ~n_13483;
assign n_13485 = ~x_873 &  n_13483;
assign n_13486 = ~n_13484 & ~n_13485;
assign n_13487 =  x_872 & ~n_13474;
assign n_13488 =  x_104 &  n_13474;
assign n_13489 = ~n_13487 & ~n_13488;
assign n_13490 =  x_872 & ~n_13489;
assign n_13491 = ~x_872 &  n_13489;
assign n_13492 = ~n_13490 & ~n_13491;
assign n_13493 =  x_871 & ~n_13474;
assign n_13494 =  x_103 &  n_13474;
assign n_13495 = ~n_13493 & ~n_13494;
assign n_13496 =  x_871 & ~n_13495;
assign n_13497 = ~x_871 &  n_13495;
assign n_13498 = ~n_13496 & ~n_13497;
assign n_13499 =  x_870 & ~n_13474;
assign n_13500 =  x_102 &  n_13474;
assign n_13501 = ~n_13499 & ~n_13500;
assign n_13502 =  x_870 & ~n_13501;
assign n_13503 = ~x_870 &  n_13501;
assign n_13504 = ~n_13502 & ~n_13503;
assign n_13505 =  x_869 & ~n_13474;
assign n_13506 =  x_101 &  n_13474;
assign n_13507 = ~n_13505 & ~n_13506;
assign n_13508 =  x_869 & ~n_13507;
assign n_13509 = ~x_869 &  n_13507;
assign n_13510 = ~n_13508 & ~n_13509;
assign n_13511 =  x_868 & ~n_13474;
assign n_13512 =  x_100 &  n_13474;
assign n_13513 = ~n_13511 & ~n_13512;
assign n_13514 =  x_868 & ~n_13513;
assign n_13515 = ~x_868 &  n_13513;
assign n_13516 = ~n_13514 & ~n_13515;
assign n_13517 =  x_867 & ~n_13474;
assign n_13518 =  x_99 &  n_13474;
assign n_13519 = ~n_13517 & ~n_13518;
assign n_13520 =  x_867 & ~n_13519;
assign n_13521 = ~x_867 &  n_13519;
assign n_13522 = ~n_13520 & ~n_13521;
assign n_13523 =  x_866 & ~n_13474;
assign n_13524 =  x_98 &  n_13474;
assign n_13525 = ~n_13523 & ~n_13524;
assign n_13526 =  x_866 & ~n_13525;
assign n_13527 = ~x_866 &  n_13525;
assign n_13528 = ~n_13526 & ~n_13527;
assign n_13529 =  x_865 & ~n_13474;
assign n_13530 =  x_97 &  n_13474;
assign n_13531 = ~n_13529 & ~n_13530;
assign n_13532 =  x_865 & ~n_13531;
assign n_13533 = ~x_865 &  n_13531;
assign n_13534 = ~n_13532 & ~n_13533;
assign n_13535 =  x_864 & ~n_13474;
assign n_13536 =  x_96 &  n_13474;
assign n_13537 = ~n_13535 & ~n_13536;
assign n_13538 =  x_864 & ~n_13537;
assign n_13539 = ~x_864 &  n_13537;
assign n_13540 = ~n_13538 & ~n_13539;
assign n_13541 =  x_863 & ~n_13474;
assign n_13542 =  x_95 &  n_13474;
assign n_13543 = ~n_13541 & ~n_13542;
assign n_13544 =  x_863 & ~n_13543;
assign n_13545 = ~x_863 &  n_13543;
assign n_13546 = ~n_13544 & ~n_13545;
assign n_13547 =  x_862 & ~n_13474;
assign n_13548 =  x_94 &  n_13474;
assign n_13549 = ~n_13547 & ~n_13548;
assign n_13550 =  x_862 & ~n_13549;
assign n_13551 = ~x_862 &  n_13549;
assign n_13552 = ~n_13550 & ~n_13551;
assign n_13553 =  x_861 & ~n_13474;
assign n_13554 =  x_93 &  n_13474;
assign n_13555 = ~n_13553 & ~n_13554;
assign n_13556 =  x_861 & ~n_13555;
assign n_13557 = ~x_861 &  n_13555;
assign n_13558 = ~n_13556 & ~n_13557;
assign n_13559 =  x_860 & ~n_13474;
assign n_13560 =  x_92 &  n_13474;
assign n_13561 = ~n_13559 & ~n_13560;
assign n_13562 =  x_860 & ~n_13561;
assign n_13563 = ~x_860 &  n_13561;
assign n_13564 = ~n_13562 & ~n_13563;
assign n_13565 =  x_859 & ~n_13474;
assign n_13566 =  x_91 &  n_13474;
assign n_13567 = ~n_13565 & ~n_13566;
assign n_13568 =  x_859 & ~n_13567;
assign n_13569 = ~x_859 &  n_13567;
assign n_13570 = ~n_13568 & ~n_13569;
assign n_13571 =  x_858 & ~n_13474;
assign n_13572 =  x_90 &  n_13474;
assign n_13573 = ~n_13571 & ~n_13572;
assign n_13574 =  x_858 & ~n_13573;
assign n_13575 = ~x_858 &  n_13573;
assign n_13576 = ~n_13574 & ~n_13575;
assign n_13577 =  x_857 & ~n_13474;
assign n_13578 =  x_89 &  n_13474;
assign n_13579 = ~n_13577 & ~n_13578;
assign n_13580 =  x_857 & ~n_13579;
assign n_13581 = ~x_857 &  n_13579;
assign n_13582 = ~n_13580 & ~n_13581;
assign n_13583 =  x_856 & ~n_13474;
assign n_13584 =  x_88 &  n_13474;
assign n_13585 = ~n_13583 & ~n_13584;
assign n_13586 =  x_856 & ~n_13585;
assign n_13587 = ~x_856 &  n_13585;
assign n_13588 = ~n_13586 & ~n_13587;
assign n_13589 =  x_855 & ~n_13474;
assign n_13590 =  x_87 &  n_13474;
assign n_13591 = ~n_13589 & ~n_13590;
assign n_13592 =  x_855 & ~n_13591;
assign n_13593 = ~x_855 &  n_13591;
assign n_13594 = ~n_13592 & ~n_13593;
assign n_13595 =  x_854 & ~n_13474;
assign n_13596 =  x_86 &  n_13474;
assign n_13597 = ~n_13595 & ~n_13596;
assign n_13598 =  x_854 & ~n_13597;
assign n_13599 = ~x_854 &  n_13597;
assign n_13600 = ~n_13598 & ~n_13599;
assign n_13601 =  x_853 & ~n_13474;
assign n_13602 =  x_85 &  n_13474;
assign n_13603 = ~n_13601 & ~n_13602;
assign n_13604 =  x_853 & ~n_13603;
assign n_13605 = ~x_853 &  n_13603;
assign n_13606 = ~n_13604 & ~n_13605;
assign n_13607 =  x_852 & ~n_13474;
assign n_13608 =  x_84 &  n_13474;
assign n_13609 = ~n_13607 & ~n_13608;
assign n_13610 =  x_852 & ~n_13609;
assign n_13611 = ~x_852 &  n_13609;
assign n_13612 = ~n_13610 & ~n_13611;
assign n_13613 =  x_851 & ~n_13474;
assign n_13614 =  x_83 &  n_13474;
assign n_13615 = ~n_13613 & ~n_13614;
assign n_13616 =  x_851 & ~n_13615;
assign n_13617 = ~x_851 &  n_13615;
assign n_13618 = ~n_13616 & ~n_13617;
assign n_13619 =  x_850 & ~n_13474;
assign n_13620 =  x_82 &  n_13474;
assign n_13621 = ~n_13619 & ~n_13620;
assign n_13622 =  x_850 & ~n_13621;
assign n_13623 = ~x_850 &  n_13621;
assign n_13624 = ~n_13622 & ~n_13623;
assign n_13625 =  x_849 & ~n_13474;
assign n_13626 =  x_81 &  n_13474;
assign n_13627 = ~n_13625 & ~n_13626;
assign n_13628 =  x_849 & ~n_13627;
assign n_13629 = ~x_849 &  n_13627;
assign n_13630 = ~n_13628 & ~n_13629;
assign n_13631 =  x_848 & ~n_13474;
assign n_13632 =  x_80 &  n_13474;
assign n_13633 = ~n_13631 & ~n_13632;
assign n_13634 =  x_848 & ~n_13633;
assign n_13635 = ~x_848 &  n_13633;
assign n_13636 = ~n_13634 & ~n_13635;
assign n_13637 =  x_847 & ~n_13474;
assign n_13638 =  x_79 &  n_13474;
assign n_13639 = ~n_13637 & ~n_13638;
assign n_13640 =  x_847 & ~n_13639;
assign n_13641 = ~x_847 &  n_13639;
assign n_13642 = ~n_13640 & ~n_13641;
assign n_13643 =  x_846 & ~n_13474;
assign n_13644 =  x_78 &  n_13474;
assign n_13645 = ~n_13643 & ~n_13644;
assign n_13646 =  x_846 & ~n_13645;
assign n_13647 = ~x_846 &  n_13645;
assign n_13648 = ~n_13646 & ~n_13647;
assign n_13649 =  x_845 & ~n_13474;
assign n_13650 =  x_77 &  n_13474;
assign n_13651 = ~n_13649 & ~n_13650;
assign n_13652 =  x_845 & ~n_13651;
assign n_13653 = ~x_845 &  n_13651;
assign n_13654 = ~n_13652 & ~n_13653;
assign n_13655 =  x_844 & ~n_13474;
assign n_13656 =  x_76 &  n_13474;
assign n_13657 = ~n_13655 & ~n_13656;
assign n_13658 =  x_844 & ~n_13657;
assign n_13659 = ~x_844 &  n_13657;
assign n_13660 = ~n_13658 & ~n_13659;
assign n_13661 =  x_843 & ~n_13474;
assign n_13662 =  x_75 &  n_13474;
assign n_13663 = ~n_13661 & ~n_13662;
assign n_13664 =  x_843 & ~n_13663;
assign n_13665 = ~x_843 &  n_13663;
assign n_13666 = ~n_13664 & ~n_13665;
assign n_13667 =  n_3 &  n_4057;
assign n_13668 =  x_842 & ~n_13667;
assign n_13669 =  i_32 &  n_13667;
assign n_13670 = ~n_13668 & ~n_13669;
assign n_13671 =  x_842 & ~n_13670;
assign n_13672 = ~x_842 &  n_13670;
assign n_13673 = ~n_13671 & ~n_13672;
assign n_13674 =  x_841 & ~n_13667;
assign n_13675 =  i_31 &  n_13667;
assign n_13676 = ~n_13674 & ~n_13675;
assign n_13677 =  x_841 & ~n_13676;
assign n_13678 = ~x_841 &  n_13676;
assign n_13679 = ~n_13677 & ~n_13678;
assign n_13680 =  x_840 & ~n_13667;
assign n_13681 =  i_30 &  n_13667;
assign n_13682 = ~n_13680 & ~n_13681;
assign n_13683 =  x_840 & ~n_13682;
assign n_13684 = ~x_840 &  n_13682;
assign n_13685 = ~n_13683 & ~n_13684;
assign n_13686 =  x_839 & ~n_13667;
assign n_13687 =  i_29 &  n_13667;
assign n_13688 = ~n_13686 & ~n_13687;
assign n_13689 =  x_839 & ~n_13688;
assign n_13690 = ~x_839 &  n_13688;
assign n_13691 = ~n_13689 & ~n_13690;
assign n_13692 =  x_838 & ~n_13667;
assign n_13693 =  i_28 &  n_13667;
assign n_13694 = ~n_13692 & ~n_13693;
assign n_13695 =  x_838 & ~n_13694;
assign n_13696 = ~x_838 &  n_13694;
assign n_13697 = ~n_13695 & ~n_13696;
assign n_13698 =  x_837 & ~n_13667;
assign n_13699 =  i_27 &  n_13667;
assign n_13700 = ~n_13698 & ~n_13699;
assign n_13701 =  x_837 & ~n_13700;
assign n_13702 = ~x_837 &  n_13700;
assign n_13703 = ~n_13701 & ~n_13702;
assign n_13704 =  x_836 & ~n_13667;
assign n_13705 =  i_26 &  n_13667;
assign n_13706 = ~n_13704 & ~n_13705;
assign n_13707 =  x_836 & ~n_13706;
assign n_13708 = ~x_836 &  n_13706;
assign n_13709 = ~n_13707 & ~n_13708;
assign n_13710 =  x_835 & ~n_13667;
assign n_13711 =  i_25 &  n_13667;
assign n_13712 = ~n_13710 & ~n_13711;
assign n_13713 =  x_835 & ~n_13712;
assign n_13714 = ~x_835 &  n_13712;
assign n_13715 = ~n_13713 & ~n_13714;
assign n_13716 =  x_834 & ~n_13667;
assign n_13717 =  i_24 &  n_13667;
assign n_13718 = ~n_13716 & ~n_13717;
assign n_13719 =  x_834 & ~n_13718;
assign n_13720 = ~x_834 &  n_13718;
assign n_13721 = ~n_13719 & ~n_13720;
assign n_13722 =  x_833 & ~n_13667;
assign n_13723 =  i_23 &  n_13667;
assign n_13724 = ~n_13722 & ~n_13723;
assign n_13725 =  x_833 & ~n_13724;
assign n_13726 = ~x_833 &  n_13724;
assign n_13727 = ~n_13725 & ~n_13726;
assign n_13728 =  x_832 & ~n_13667;
assign n_13729 =  i_22 &  n_13667;
assign n_13730 = ~n_13728 & ~n_13729;
assign n_13731 =  x_832 & ~n_13730;
assign n_13732 = ~x_832 &  n_13730;
assign n_13733 = ~n_13731 & ~n_13732;
assign n_13734 =  x_831 & ~n_13667;
assign n_13735 =  i_21 &  n_13667;
assign n_13736 = ~n_13734 & ~n_13735;
assign n_13737 =  x_831 & ~n_13736;
assign n_13738 = ~x_831 &  n_13736;
assign n_13739 = ~n_13737 & ~n_13738;
assign n_13740 =  x_830 & ~n_13667;
assign n_13741 =  i_20 &  n_13667;
assign n_13742 = ~n_13740 & ~n_13741;
assign n_13743 =  x_830 & ~n_13742;
assign n_13744 = ~x_830 &  n_13742;
assign n_13745 = ~n_13743 & ~n_13744;
assign n_13746 =  x_829 & ~n_13667;
assign n_13747 =  i_19 &  n_13667;
assign n_13748 = ~n_13746 & ~n_13747;
assign n_13749 =  x_829 & ~n_13748;
assign n_13750 = ~x_829 &  n_13748;
assign n_13751 = ~n_13749 & ~n_13750;
assign n_13752 =  x_828 & ~n_13667;
assign n_13753 =  i_18 &  n_13667;
assign n_13754 = ~n_13752 & ~n_13753;
assign n_13755 =  x_828 & ~n_13754;
assign n_13756 = ~x_828 &  n_13754;
assign n_13757 = ~n_13755 & ~n_13756;
assign n_13758 =  x_827 & ~n_13667;
assign n_13759 =  i_17 &  n_13667;
assign n_13760 = ~n_13758 & ~n_13759;
assign n_13761 =  x_827 & ~n_13760;
assign n_13762 = ~x_827 &  n_13760;
assign n_13763 = ~n_13761 & ~n_13762;
assign n_13764 =  x_826 & ~n_13667;
assign n_13765 =  i_16 &  n_13667;
assign n_13766 = ~n_13764 & ~n_13765;
assign n_13767 =  x_826 & ~n_13766;
assign n_13768 = ~x_826 &  n_13766;
assign n_13769 = ~n_13767 & ~n_13768;
assign n_13770 =  x_825 & ~n_13667;
assign n_13771 =  i_15 &  n_13667;
assign n_13772 = ~n_13770 & ~n_13771;
assign n_13773 =  x_825 & ~n_13772;
assign n_13774 = ~x_825 &  n_13772;
assign n_13775 = ~n_13773 & ~n_13774;
assign n_13776 =  x_824 & ~n_13667;
assign n_13777 =  i_14 &  n_13667;
assign n_13778 = ~n_13776 & ~n_13777;
assign n_13779 =  x_824 & ~n_13778;
assign n_13780 = ~x_824 &  n_13778;
assign n_13781 = ~n_13779 & ~n_13780;
assign n_13782 =  x_823 & ~n_13667;
assign n_13783 =  i_13 &  n_13667;
assign n_13784 = ~n_13782 & ~n_13783;
assign n_13785 =  x_823 & ~n_13784;
assign n_13786 = ~x_823 &  n_13784;
assign n_13787 = ~n_13785 & ~n_13786;
assign n_13788 =  x_822 & ~n_13667;
assign n_13789 =  i_12 &  n_13667;
assign n_13790 = ~n_13788 & ~n_13789;
assign n_13791 =  x_822 & ~n_13790;
assign n_13792 = ~x_822 &  n_13790;
assign n_13793 = ~n_13791 & ~n_13792;
assign n_13794 =  x_821 & ~n_13667;
assign n_13795 =  i_11 &  n_13667;
assign n_13796 = ~n_13794 & ~n_13795;
assign n_13797 =  x_821 & ~n_13796;
assign n_13798 = ~x_821 &  n_13796;
assign n_13799 = ~n_13797 & ~n_13798;
assign n_13800 =  x_820 & ~n_13667;
assign n_13801 =  i_10 &  n_13667;
assign n_13802 = ~n_13800 & ~n_13801;
assign n_13803 =  x_820 & ~n_13802;
assign n_13804 = ~x_820 &  n_13802;
assign n_13805 = ~n_13803 & ~n_13804;
assign n_13806 =  x_819 & ~n_13667;
assign n_13807 =  i_9 &  n_13667;
assign n_13808 = ~n_13806 & ~n_13807;
assign n_13809 =  x_819 & ~n_13808;
assign n_13810 = ~x_819 &  n_13808;
assign n_13811 = ~n_13809 & ~n_13810;
assign n_13812 =  x_818 & ~n_13667;
assign n_13813 =  i_8 &  n_13667;
assign n_13814 = ~n_13812 & ~n_13813;
assign n_13815 =  x_818 & ~n_13814;
assign n_13816 = ~x_818 &  n_13814;
assign n_13817 = ~n_13815 & ~n_13816;
assign n_13818 =  x_817 & ~n_13667;
assign n_13819 =  i_7 &  n_13667;
assign n_13820 = ~n_13818 & ~n_13819;
assign n_13821 =  x_817 & ~n_13820;
assign n_13822 = ~x_817 &  n_13820;
assign n_13823 = ~n_13821 & ~n_13822;
assign n_13824 =  x_816 & ~n_13667;
assign n_13825 =  i_6 &  n_13667;
assign n_13826 = ~n_13824 & ~n_13825;
assign n_13827 =  x_816 & ~n_13826;
assign n_13828 = ~x_816 &  n_13826;
assign n_13829 = ~n_13827 & ~n_13828;
assign n_13830 =  x_815 & ~n_13667;
assign n_13831 =  i_5 &  n_13667;
assign n_13832 = ~n_13830 & ~n_13831;
assign n_13833 =  x_815 & ~n_13832;
assign n_13834 = ~x_815 &  n_13832;
assign n_13835 = ~n_13833 & ~n_13834;
assign n_13836 =  x_814 & ~n_13667;
assign n_13837 =  i_4 &  n_13667;
assign n_13838 = ~n_13836 & ~n_13837;
assign n_13839 =  x_814 & ~n_13838;
assign n_13840 = ~x_814 &  n_13838;
assign n_13841 = ~n_13839 & ~n_13840;
assign n_13842 =  x_813 & ~n_13667;
assign n_13843 =  i_3 &  n_13667;
assign n_13844 = ~n_13842 & ~n_13843;
assign n_13845 =  x_813 & ~n_13844;
assign n_13846 = ~x_813 &  n_13844;
assign n_13847 = ~n_13845 & ~n_13846;
assign n_13848 =  x_812 & ~n_13667;
assign n_13849 =  i_2 &  n_13667;
assign n_13850 = ~n_13848 & ~n_13849;
assign n_13851 =  x_812 & ~n_13850;
assign n_13852 = ~x_812 &  n_13850;
assign n_13853 = ~n_13851 & ~n_13852;
assign n_13854 =  x_811 & ~n_13667;
assign n_13855 =  i_1 &  n_13667;
assign n_13856 = ~n_13854 & ~n_13855;
assign n_13857 =  x_811 & ~n_13856;
assign n_13858 = ~x_811 &  n_13856;
assign n_13859 = ~n_13857 & ~n_13858;
assign n_13860 =  x_41 &  n_391;
assign n_13861 =  x_2314 &  x_2730;
assign n_13862 = ~x_2314 & ~x_2730;
assign n_13863 = ~n_13861 & ~n_13862;
assign n_13864 =  n_13860 &  n_13863;
assign n_13865 =  n_3858 & ~n_3861;
assign n_13866 =  n_3860 &  n_13865;
assign n_13867 =  x_810 & ~n_13866;
assign n_13868 =  n_184 &  n_390;
assign n_13869 =  n_185 &  n_13868;
assign n_13870 =  x_490 &  x_1226;
assign n_13871 = ~x_490 & ~x_1226;
assign n_13872 = ~n_13870 & ~n_13871;
assign n_13873 =  n_13869 &  n_13872;
assign n_13874 = ~n_13867 & ~n_13873;
assign n_13875 = ~n_13864 &  n_13874;
assign n_13876 =  x_810 & ~n_13875;
assign n_13877 = ~x_810 &  n_13875;
assign n_13878 = ~n_13876 & ~n_13877;
assign n_13879 = ~x_489 & ~x_490;
assign n_13880 =  x_489 &  x_490;
assign n_13881 = ~n_13879 & ~n_13880;
assign n_13882 =  x_1225 &  n_13881;
assign n_13883 = ~x_1225 & ~n_13881;
assign n_13884 = ~n_13882 & ~n_13883;
assign n_13885 =  n_13870 &  n_13884;
assign n_13886 = ~n_13870 & ~n_13884;
assign n_13887 = ~n_13885 & ~n_13886;
assign n_13888 =  n_13869 &  n_13887;
assign n_13889 =  x_809 & ~n_13866;
assign n_13890 = ~x_2729 & ~x_2730;
assign n_13891 =  x_2729 &  x_2730;
assign n_13892 = ~n_13890 & ~n_13891;
assign n_13893 =  x_2313 &  n_13892;
assign n_13894 = ~x_2313 & ~n_13892;
assign n_13895 = ~n_13893 & ~n_13894;
assign n_13896 =  n_13861 &  n_13895;
assign n_13897 = ~n_13861 & ~n_13895;
assign n_13898 = ~n_13896 & ~n_13897;
assign n_13899 =  n_13860 &  n_13898;
assign n_13900 = ~n_13889 & ~n_13899;
assign n_13901 = ~n_13888 &  n_13900;
assign n_13902 =  x_809 & ~n_13901;
assign n_13903 = ~x_809 &  n_13901;
assign n_13904 = ~n_13902 & ~n_13903;
assign n_13905 = ~x_488 &  n_13879;
assign n_13906 =  x_488 & ~n_13879;
assign n_13907 = ~n_13905 & ~n_13906;
assign n_13908 =  x_489 & ~x_1225;
assign n_13909 =  n_13870 & ~n_13908;
assign n_13910 = ~n_13909 & ~n_13882;
assign n_13911 =  n_13907 & ~n_13910;
assign n_13912 = ~n_13907 &  n_13910;
assign n_13913 = ~n_13911 & ~n_13912;
assign n_13914 = ~x_1224 & ~n_13913;
assign n_13915 =  x_1224 & ~n_13912;
assign n_13916 = ~n_13911 &  n_13915;
assign n_13917 =  n_13869 & ~n_13916;
assign n_13918 = ~n_13914 &  n_13917;
assign n_13919 =  x_808 & ~n_13866;
assign n_13920 = ~x_2728 &  n_13890;
assign n_13921 =  x_2728 & ~n_13890;
assign n_13922 = ~n_13920 & ~n_13921;
assign n_13923 = ~x_2313 &  x_2729;
assign n_13924 =  n_13861 & ~n_13923;
assign n_13925 = ~n_13924 & ~n_13893;
assign n_13926 =  n_13922 & ~n_13925;
assign n_13927 = ~n_13922 &  n_13925;
assign n_13928 = ~n_13926 & ~n_13927;
assign n_13929 = ~x_2312 & ~n_13928;
assign n_13930 =  x_2312 & ~n_13927;
assign n_13931 = ~n_13926 &  n_13930;
assign n_13932 =  n_13860 & ~n_13931;
assign n_13933 = ~n_13929 &  n_13932;
assign n_13934 = ~n_13919 & ~n_13933;
assign n_13935 = ~n_13918 &  n_13934;
assign n_13936 =  x_808 & ~n_13935;
assign n_13937 = ~x_808 &  n_13935;
assign n_13938 = ~n_13936 & ~n_13937;
assign n_13939 = ~x_2727 &  n_13920;
assign n_13940 =  x_2727 & ~n_13920;
assign n_13941 = ~n_13939 & ~n_13940;
assign n_13942 = ~n_13926 & ~n_13930;
assign n_13943 =  n_13941 & ~n_13942;
assign n_13944 = ~n_13941 &  n_13942;
assign n_13945 = ~n_13943 & ~n_13944;
assign n_13946 = ~x_2311 & ~n_13945;
assign n_13947 =  x_2311 & ~n_13944;
assign n_13948 = ~n_13943 &  n_13947;
assign n_13949 =  n_13860 & ~n_13948;
assign n_13950 = ~n_13946 &  n_13949;
assign n_13951 =  x_807 & ~n_13866;
assign n_13952 = ~x_487 &  n_13905;
assign n_13953 =  x_487 & ~n_13905;
assign n_13954 = ~n_13952 & ~n_13953;
assign n_13955 = ~n_13911 & ~n_13915;
assign n_13956 =  n_13954 & ~n_13955;
assign n_13957 = ~n_13954 &  n_13955;
assign n_13958 = ~n_13956 & ~n_13957;
assign n_13959 = ~x_1223 & ~n_13958;
assign n_13960 =  x_1223 & ~n_13957;
assign n_13961 = ~n_13956 &  n_13960;
assign n_13962 =  n_13869 & ~n_13961;
assign n_13963 = ~n_13959 &  n_13962;
assign n_13964 = ~n_13951 & ~n_13963;
assign n_13965 = ~n_13950 &  n_13964;
assign n_13966 =  x_807 & ~n_13965;
assign n_13967 = ~x_807 &  n_13965;
assign n_13968 = ~n_13966 & ~n_13967;
assign n_13969 = ~x_2726 &  n_13939;
assign n_13970 =  x_2726 & ~n_13939;
assign n_13971 = ~n_13969 & ~n_13970;
assign n_13972 = ~n_13943 & ~n_13947;
assign n_13973 =  n_13971 & ~n_13972;
assign n_13974 = ~n_13971 &  n_13972;
assign n_13975 = ~n_13973 & ~n_13974;
assign n_13976 = ~x_2310 & ~n_13975;
assign n_13977 =  x_2310 & ~n_13974;
assign n_13978 = ~n_13973 &  n_13977;
assign n_13979 =  n_13860 & ~n_13978;
assign n_13980 = ~n_13976 &  n_13979;
assign n_13981 =  x_806 & ~n_13866;
assign n_13982 = ~x_486 &  n_13952;
assign n_13983 =  x_486 & ~n_13952;
assign n_13984 = ~n_13982 & ~n_13983;
assign n_13985 = ~n_13956 & ~n_13960;
assign n_13986 =  n_13984 & ~n_13985;
assign n_13987 = ~n_13984 &  n_13985;
assign n_13988 = ~n_13986 & ~n_13987;
assign n_13989 = ~x_1222 & ~n_13988;
assign n_13990 =  x_1222 & ~n_13987;
assign n_13991 = ~n_13986 &  n_13990;
assign n_13992 =  n_13869 & ~n_13991;
assign n_13993 = ~n_13989 &  n_13992;
assign n_13994 = ~n_13981 & ~n_13993;
assign n_13995 = ~n_13980 &  n_13994;
assign n_13996 =  x_806 & ~n_13995;
assign n_13997 = ~x_806 &  n_13995;
assign n_13998 = ~n_13996 & ~n_13997;
assign n_13999 = ~x_2725 &  n_13969;
assign n_14000 =  x_2725 & ~n_13969;
assign n_14001 = ~n_13999 & ~n_14000;
assign n_14002 = ~n_13973 & ~n_13977;
assign n_14003 =  n_14001 & ~n_14002;
assign n_14004 = ~n_14001 &  n_14002;
assign n_14005 = ~n_14003 & ~n_14004;
assign n_14006 = ~x_2309 & ~n_14005;
assign n_14007 =  x_2309 & ~n_14004;
assign n_14008 = ~n_14003 &  n_14007;
assign n_14009 =  n_13860 & ~n_14008;
assign n_14010 = ~n_14006 &  n_14009;
assign n_14011 =  x_805 & ~n_13866;
assign n_14012 = ~x_485 &  n_13982;
assign n_14013 =  x_485 & ~n_13982;
assign n_14014 = ~n_14012 & ~n_14013;
assign n_14015 = ~n_13986 & ~n_13990;
assign n_14016 =  n_14014 & ~n_14015;
assign n_14017 = ~n_14014 &  n_14015;
assign n_14018 = ~n_14016 & ~n_14017;
assign n_14019 = ~x_1221 & ~n_14018;
assign n_14020 =  x_1221 & ~n_14017;
assign n_14021 = ~n_14016 &  n_14020;
assign n_14022 =  n_13869 & ~n_14021;
assign n_14023 = ~n_14019 &  n_14022;
assign n_14024 = ~n_14011 & ~n_14023;
assign n_14025 = ~n_14010 &  n_14024;
assign n_14026 =  x_805 & ~n_14025;
assign n_14027 = ~x_805 &  n_14025;
assign n_14028 = ~n_14026 & ~n_14027;
assign n_14029 = ~x_2724 &  n_13999;
assign n_14030 =  x_2724 & ~n_13999;
assign n_14031 = ~n_14029 & ~n_14030;
assign n_14032 = ~n_14003 & ~n_14007;
assign n_14033 =  n_14031 & ~n_14032;
assign n_14034 = ~n_14031 &  n_14032;
assign n_14035 = ~n_14033 & ~n_14034;
assign n_14036 = ~x_2308 & ~n_14035;
assign n_14037 =  x_2308 & ~n_14034;
assign n_14038 = ~n_14033 &  n_14037;
assign n_14039 =  n_13860 & ~n_14038;
assign n_14040 = ~n_14036 &  n_14039;
assign n_14041 =  x_804 & ~n_13866;
assign n_14042 = ~x_484 &  n_14012;
assign n_14043 =  x_484 & ~n_14012;
assign n_14044 = ~n_14042 & ~n_14043;
assign n_14045 = ~n_14016 & ~n_14020;
assign n_14046 =  n_14044 & ~n_14045;
assign n_14047 = ~n_14044 &  n_14045;
assign n_14048 = ~n_14046 & ~n_14047;
assign n_14049 = ~x_1220 & ~n_14048;
assign n_14050 =  x_1220 & ~n_14047;
assign n_14051 = ~n_14046 &  n_14050;
assign n_14052 =  n_13869 & ~n_14051;
assign n_14053 = ~n_14049 &  n_14052;
assign n_14054 = ~n_14041 & ~n_14053;
assign n_14055 = ~n_14040 &  n_14054;
assign n_14056 =  x_804 & ~n_14055;
assign n_14057 = ~x_804 &  n_14055;
assign n_14058 = ~n_14056 & ~n_14057;
assign n_14059 = ~x_2723 &  n_14029;
assign n_14060 =  x_2723 & ~n_14029;
assign n_14061 = ~n_14059 & ~n_14060;
assign n_14062 = ~n_14033 & ~n_14037;
assign n_14063 =  n_14061 & ~n_14062;
assign n_14064 = ~n_14061 &  n_14062;
assign n_14065 = ~n_14063 & ~n_14064;
assign n_14066 = ~x_2307 & ~n_14065;
assign n_14067 =  x_2307 & ~n_14064;
assign n_14068 = ~n_14063 &  n_14067;
assign n_14069 =  n_13860 & ~n_14068;
assign n_14070 = ~n_14066 &  n_14069;
assign n_14071 =  x_803 & ~n_13866;
assign n_14072 = ~x_483 &  n_14042;
assign n_14073 =  x_483 & ~n_14042;
assign n_14074 = ~n_14072 & ~n_14073;
assign n_14075 = ~n_14046 & ~n_14050;
assign n_14076 =  n_14074 & ~n_14075;
assign n_14077 = ~n_14074 &  n_14075;
assign n_14078 = ~n_14076 & ~n_14077;
assign n_14079 = ~x_1219 & ~n_14078;
assign n_14080 =  x_1219 & ~n_14077;
assign n_14081 = ~n_14076 &  n_14080;
assign n_14082 =  n_13869 & ~n_14081;
assign n_14083 = ~n_14079 &  n_14082;
assign n_14084 = ~n_14071 & ~n_14083;
assign n_14085 = ~n_14070 &  n_14084;
assign n_14086 =  x_803 & ~n_14085;
assign n_14087 = ~x_803 &  n_14085;
assign n_14088 = ~n_14086 & ~n_14087;
assign n_14089 = ~x_2722 &  n_14059;
assign n_14090 =  x_2722 & ~n_14059;
assign n_14091 = ~n_14089 & ~n_14090;
assign n_14092 = ~n_14063 & ~n_14067;
assign n_14093 =  n_14091 & ~n_14092;
assign n_14094 = ~n_14091 &  n_14092;
assign n_14095 = ~n_14093 & ~n_14094;
assign n_14096 = ~x_2306 & ~n_14095;
assign n_14097 =  x_2306 & ~n_14094;
assign n_14098 = ~n_14093 &  n_14097;
assign n_14099 =  n_13860 & ~n_14098;
assign n_14100 = ~n_14096 &  n_14099;
assign n_14101 =  x_802 & ~n_13866;
assign n_14102 = ~x_482 &  n_14072;
assign n_14103 =  x_482 & ~n_14072;
assign n_14104 = ~n_14102 & ~n_14103;
assign n_14105 = ~n_14076 & ~n_14080;
assign n_14106 =  n_14104 & ~n_14105;
assign n_14107 = ~n_14104 &  n_14105;
assign n_14108 = ~n_14106 & ~n_14107;
assign n_14109 = ~x_1218 & ~n_14108;
assign n_14110 =  x_1218 & ~n_14107;
assign n_14111 = ~n_14106 &  n_14110;
assign n_14112 =  n_13869 & ~n_14111;
assign n_14113 = ~n_14109 &  n_14112;
assign n_14114 = ~n_14101 & ~n_14113;
assign n_14115 = ~n_14100 &  n_14114;
assign n_14116 =  x_802 & ~n_14115;
assign n_14117 = ~x_802 &  n_14115;
assign n_14118 = ~n_14116 & ~n_14117;
assign n_14119 = ~x_2721 &  n_14089;
assign n_14120 =  x_2721 & ~n_14089;
assign n_14121 = ~n_14119 & ~n_14120;
assign n_14122 = ~n_14093 & ~n_14097;
assign n_14123 =  n_14121 & ~n_14122;
assign n_14124 = ~n_14121 &  n_14122;
assign n_14125 = ~n_14123 & ~n_14124;
assign n_14126 = ~x_2305 & ~n_14125;
assign n_14127 =  x_2305 & ~n_14124;
assign n_14128 = ~n_14123 &  n_14127;
assign n_14129 =  n_13860 & ~n_14128;
assign n_14130 = ~n_14126 &  n_14129;
assign n_14131 =  x_801 & ~n_13866;
assign n_14132 = ~x_481 &  n_14102;
assign n_14133 =  x_481 & ~n_14102;
assign n_14134 = ~n_14132 & ~n_14133;
assign n_14135 = ~n_14106 & ~n_14110;
assign n_14136 =  n_14134 & ~n_14135;
assign n_14137 = ~n_14134 &  n_14135;
assign n_14138 = ~n_14136 & ~n_14137;
assign n_14139 = ~x_1217 & ~n_14138;
assign n_14140 =  x_1217 & ~n_14137;
assign n_14141 = ~n_14136 &  n_14140;
assign n_14142 =  n_13869 & ~n_14141;
assign n_14143 = ~n_14139 &  n_14142;
assign n_14144 = ~n_14131 & ~n_14143;
assign n_14145 = ~n_14130 &  n_14144;
assign n_14146 =  x_801 & ~n_14145;
assign n_14147 = ~x_801 &  n_14145;
assign n_14148 = ~n_14146 & ~n_14147;
assign n_14149 = ~x_2720 &  n_14119;
assign n_14150 =  x_2720 & ~n_14119;
assign n_14151 = ~n_14149 & ~n_14150;
assign n_14152 = ~n_14123 & ~n_14127;
assign n_14153 =  n_14151 & ~n_14152;
assign n_14154 = ~n_14151 &  n_14152;
assign n_14155 = ~n_14153 & ~n_14154;
assign n_14156 = ~x_2304 & ~n_14155;
assign n_14157 =  x_2304 & ~n_14154;
assign n_14158 = ~n_14153 &  n_14157;
assign n_14159 =  n_13860 & ~n_14158;
assign n_14160 = ~n_14156 &  n_14159;
assign n_14161 =  x_800 & ~n_13866;
assign n_14162 = ~x_480 &  n_14132;
assign n_14163 =  x_480 & ~n_14132;
assign n_14164 = ~n_14162 & ~n_14163;
assign n_14165 = ~n_14136 & ~n_14140;
assign n_14166 =  n_14164 & ~n_14165;
assign n_14167 = ~n_14164 &  n_14165;
assign n_14168 = ~n_14166 & ~n_14167;
assign n_14169 = ~x_1216 & ~n_14168;
assign n_14170 =  x_1216 & ~n_14167;
assign n_14171 = ~n_14166 &  n_14170;
assign n_14172 =  n_13869 & ~n_14171;
assign n_14173 = ~n_14169 &  n_14172;
assign n_14174 = ~n_14161 & ~n_14173;
assign n_14175 = ~n_14160 &  n_14174;
assign n_14176 =  x_800 & ~n_14175;
assign n_14177 = ~x_800 &  n_14175;
assign n_14178 = ~n_14176 & ~n_14177;
assign n_14179 = ~x_2719 &  n_14149;
assign n_14180 =  x_2719 & ~n_14149;
assign n_14181 = ~n_14179 & ~n_14180;
assign n_14182 = ~n_14153 & ~n_14157;
assign n_14183 =  n_14181 & ~n_14182;
assign n_14184 = ~n_14181 &  n_14182;
assign n_14185 = ~n_14183 & ~n_14184;
assign n_14186 = ~x_2303 & ~n_14185;
assign n_14187 =  x_2303 & ~n_14184;
assign n_14188 = ~n_14183 &  n_14187;
assign n_14189 =  n_13860 & ~n_14188;
assign n_14190 = ~n_14186 &  n_14189;
assign n_14191 =  x_799 & ~n_13866;
assign n_14192 = ~x_479 &  n_14162;
assign n_14193 =  x_479 & ~n_14162;
assign n_14194 = ~n_14192 & ~n_14193;
assign n_14195 = ~n_14166 & ~n_14170;
assign n_14196 =  n_14194 & ~n_14195;
assign n_14197 = ~n_14194 &  n_14195;
assign n_14198 = ~n_14196 & ~n_14197;
assign n_14199 = ~x_1215 & ~n_14198;
assign n_14200 =  x_1215 & ~n_14197;
assign n_14201 = ~n_14196 &  n_14200;
assign n_14202 =  n_13869 & ~n_14201;
assign n_14203 = ~n_14199 &  n_14202;
assign n_14204 = ~n_14191 & ~n_14203;
assign n_14205 = ~n_14190 &  n_14204;
assign n_14206 =  x_799 & ~n_14205;
assign n_14207 = ~x_799 &  n_14205;
assign n_14208 = ~n_14206 & ~n_14207;
assign n_14209 = ~x_2718 &  n_14179;
assign n_14210 =  x_2718 & ~n_14179;
assign n_14211 = ~n_14209 & ~n_14210;
assign n_14212 = ~n_14183 & ~n_14187;
assign n_14213 =  n_14211 & ~n_14212;
assign n_14214 = ~n_14211 &  n_14212;
assign n_14215 = ~n_14213 & ~n_14214;
assign n_14216 = ~x_2302 & ~n_14215;
assign n_14217 =  x_2302 & ~n_14214;
assign n_14218 = ~n_14213 &  n_14217;
assign n_14219 =  n_13860 & ~n_14218;
assign n_14220 = ~n_14216 &  n_14219;
assign n_14221 =  x_798 & ~n_13866;
assign n_14222 = ~x_478 &  n_14192;
assign n_14223 =  x_478 & ~n_14192;
assign n_14224 = ~n_14222 & ~n_14223;
assign n_14225 = ~n_14196 & ~n_14200;
assign n_14226 =  n_14224 & ~n_14225;
assign n_14227 = ~n_14224 &  n_14225;
assign n_14228 = ~n_14226 & ~n_14227;
assign n_14229 = ~x_1214 & ~n_14228;
assign n_14230 =  x_1214 & ~n_14227;
assign n_14231 = ~n_14226 &  n_14230;
assign n_14232 =  n_13869 & ~n_14231;
assign n_14233 = ~n_14229 &  n_14232;
assign n_14234 = ~n_14221 & ~n_14233;
assign n_14235 = ~n_14220 &  n_14234;
assign n_14236 =  x_798 & ~n_14235;
assign n_14237 = ~x_798 &  n_14235;
assign n_14238 = ~n_14236 & ~n_14237;
assign n_14239 = ~x_2717 &  n_14209;
assign n_14240 =  x_2717 & ~n_14209;
assign n_14241 = ~n_14239 & ~n_14240;
assign n_14242 = ~n_14213 & ~n_14217;
assign n_14243 =  n_14241 & ~n_14242;
assign n_14244 = ~n_14241 &  n_14242;
assign n_14245 = ~n_14243 & ~n_14244;
assign n_14246 = ~x_2301 & ~n_14245;
assign n_14247 =  x_2301 & ~n_14244;
assign n_14248 = ~n_14243 &  n_14247;
assign n_14249 =  n_13860 & ~n_14248;
assign n_14250 = ~n_14246 &  n_14249;
assign n_14251 =  x_797 & ~n_13866;
assign n_14252 = ~x_477 &  n_14222;
assign n_14253 =  x_477 & ~n_14222;
assign n_14254 = ~n_14252 & ~n_14253;
assign n_14255 = ~n_14226 & ~n_14230;
assign n_14256 =  n_14254 & ~n_14255;
assign n_14257 = ~n_14254 &  n_14255;
assign n_14258 = ~n_14256 & ~n_14257;
assign n_14259 = ~x_1213 & ~n_14258;
assign n_14260 =  x_1213 & ~n_14257;
assign n_14261 = ~n_14256 &  n_14260;
assign n_14262 =  n_13869 & ~n_14261;
assign n_14263 = ~n_14259 &  n_14262;
assign n_14264 = ~n_14251 & ~n_14263;
assign n_14265 = ~n_14250 &  n_14264;
assign n_14266 =  x_797 & ~n_14265;
assign n_14267 = ~x_797 &  n_14265;
assign n_14268 = ~n_14266 & ~n_14267;
assign n_14269 = ~x_2716 &  n_14239;
assign n_14270 =  x_2716 & ~n_14239;
assign n_14271 = ~n_14269 & ~n_14270;
assign n_14272 = ~n_14243 & ~n_14247;
assign n_14273 =  n_14271 & ~n_14272;
assign n_14274 = ~n_14271 &  n_14272;
assign n_14275 = ~n_14273 & ~n_14274;
assign n_14276 = ~x_2300 & ~n_14275;
assign n_14277 =  x_2300 & ~n_14274;
assign n_14278 = ~n_14273 &  n_14277;
assign n_14279 =  n_13860 & ~n_14278;
assign n_14280 = ~n_14276 &  n_14279;
assign n_14281 =  x_796 & ~n_13866;
assign n_14282 = ~x_476 &  n_14252;
assign n_14283 =  x_476 & ~n_14252;
assign n_14284 = ~n_14282 & ~n_14283;
assign n_14285 = ~n_14256 & ~n_14260;
assign n_14286 =  n_14284 & ~n_14285;
assign n_14287 = ~n_14284 &  n_14285;
assign n_14288 = ~n_14286 & ~n_14287;
assign n_14289 = ~x_1212 & ~n_14288;
assign n_14290 =  x_1212 & ~n_14287;
assign n_14291 = ~n_14286 &  n_14290;
assign n_14292 =  n_13869 & ~n_14291;
assign n_14293 = ~n_14289 &  n_14292;
assign n_14294 = ~n_14281 & ~n_14293;
assign n_14295 = ~n_14280 &  n_14294;
assign n_14296 =  x_796 & ~n_14295;
assign n_14297 = ~x_796 &  n_14295;
assign n_14298 = ~n_14296 & ~n_14297;
assign n_14299 = ~x_2715 &  n_14269;
assign n_14300 =  x_2715 & ~n_14269;
assign n_14301 = ~n_14299 & ~n_14300;
assign n_14302 = ~n_14273 & ~n_14277;
assign n_14303 =  n_14301 & ~n_14302;
assign n_14304 = ~n_14301 &  n_14302;
assign n_14305 = ~n_14303 & ~n_14304;
assign n_14306 = ~x_2299 & ~n_14305;
assign n_14307 =  x_2299 & ~n_14304;
assign n_14308 = ~n_14303 &  n_14307;
assign n_14309 =  n_13860 & ~n_14308;
assign n_14310 = ~n_14306 &  n_14309;
assign n_14311 =  x_795 & ~n_13866;
assign n_14312 = ~x_475 &  n_14282;
assign n_14313 =  x_475 & ~n_14282;
assign n_14314 = ~n_14312 & ~n_14313;
assign n_14315 = ~n_14286 & ~n_14290;
assign n_14316 =  n_14314 & ~n_14315;
assign n_14317 = ~n_14314 &  n_14315;
assign n_14318 = ~n_14316 & ~n_14317;
assign n_14319 = ~x_1211 & ~n_14318;
assign n_14320 =  x_1211 & ~n_14317;
assign n_14321 = ~n_14316 &  n_14320;
assign n_14322 =  n_13869 & ~n_14321;
assign n_14323 = ~n_14319 &  n_14322;
assign n_14324 = ~n_14311 & ~n_14323;
assign n_14325 = ~n_14310 &  n_14324;
assign n_14326 =  x_795 & ~n_14325;
assign n_14327 = ~x_795 &  n_14325;
assign n_14328 = ~n_14326 & ~n_14327;
assign n_14329 = ~x_2714 &  n_14299;
assign n_14330 =  x_2714 & ~n_14299;
assign n_14331 = ~n_14329 & ~n_14330;
assign n_14332 = ~n_14303 & ~n_14307;
assign n_14333 =  n_14331 & ~n_14332;
assign n_14334 = ~n_14331 &  n_14332;
assign n_14335 = ~n_14333 & ~n_14334;
assign n_14336 = ~x_2298 & ~n_14335;
assign n_14337 =  x_2298 & ~n_14334;
assign n_14338 = ~n_14333 &  n_14337;
assign n_14339 =  n_13860 & ~n_14338;
assign n_14340 = ~n_14336 &  n_14339;
assign n_14341 =  x_794 & ~n_13866;
assign n_14342 = ~x_474 &  n_14312;
assign n_14343 =  x_474 & ~n_14312;
assign n_14344 = ~n_14342 & ~n_14343;
assign n_14345 = ~n_14316 & ~n_14320;
assign n_14346 =  n_14344 & ~n_14345;
assign n_14347 = ~n_14344 &  n_14345;
assign n_14348 = ~n_14346 & ~n_14347;
assign n_14349 = ~x_1210 & ~n_14348;
assign n_14350 =  x_1210 & ~n_14347;
assign n_14351 = ~n_14346 &  n_14350;
assign n_14352 =  n_13869 & ~n_14351;
assign n_14353 = ~n_14349 &  n_14352;
assign n_14354 = ~n_14341 & ~n_14353;
assign n_14355 = ~n_14340 &  n_14354;
assign n_14356 =  x_794 & ~n_14355;
assign n_14357 = ~x_794 &  n_14355;
assign n_14358 = ~n_14356 & ~n_14357;
assign n_14359 = ~x_2713 &  n_14329;
assign n_14360 =  x_2713 & ~n_14329;
assign n_14361 = ~n_14359 & ~n_14360;
assign n_14362 = ~n_14333 & ~n_14337;
assign n_14363 =  n_14361 & ~n_14362;
assign n_14364 = ~n_14361 &  n_14362;
assign n_14365 = ~n_14363 & ~n_14364;
assign n_14366 = ~x_2297 & ~n_14365;
assign n_14367 =  x_2297 & ~n_14364;
assign n_14368 = ~n_14363 &  n_14367;
assign n_14369 =  n_13860 & ~n_14368;
assign n_14370 = ~n_14366 &  n_14369;
assign n_14371 =  x_793 & ~n_13866;
assign n_14372 = ~x_473 &  n_14342;
assign n_14373 =  x_473 & ~n_14342;
assign n_14374 = ~n_14372 & ~n_14373;
assign n_14375 = ~n_14346 & ~n_14350;
assign n_14376 =  n_14374 & ~n_14375;
assign n_14377 = ~n_14374 &  n_14375;
assign n_14378 = ~n_14376 & ~n_14377;
assign n_14379 = ~x_1209 & ~n_14378;
assign n_14380 =  x_1209 & ~n_14377;
assign n_14381 = ~n_14376 &  n_14380;
assign n_14382 =  n_13869 & ~n_14381;
assign n_14383 = ~n_14379 &  n_14382;
assign n_14384 = ~n_14371 & ~n_14383;
assign n_14385 = ~n_14370 &  n_14384;
assign n_14386 =  x_793 & ~n_14385;
assign n_14387 = ~x_793 &  n_14385;
assign n_14388 = ~n_14386 & ~n_14387;
assign n_14389 = ~x_2712 &  n_14359;
assign n_14390 =  x_2712 & ~n_14359;
assign n_14391 = ~n_14389 & ~n_14390;
assign n_14392 = ~n_14363 & ~n_14367;
assign n_14393 =  n_14391 & ~n_14392;
assign n_14394 = ~n_14391 &  n_14392;
assign n_14395 = ~n_14393 & ~n_14394;
assign n_14396 = ~x_2296 & ~n_14395;
assign n_14397 =  x_2296 & ~n_14394;
assign n_14398 = ~n_14393 &  n_14397;
assign n_14399 =  n_13860 & ~n_14398;
assign n_14400 = ~n_14396 &  n_14399;
assign n_14401 =  x_792 & ~n_13866;
assign n_14402 = ~x_472 &  n_14372;
assign n_14403 =  x_472 & ~n_14372;
assign n_14404 = ~n_14402 & ~n_14403;
assign n_14405 = ~n_14376 & ~n_14380;
assign n_14406 =  n_14404 & ~n_14405;
assign n_14407 = ~n_14404 &  n_14405;
assign n_14408 = ~n_14406 & ~n_14407;
assign n_14409 = ~x_1208 & ~n_14408;
assign n_14410 =  x_1208 & ~n_14407;
assign n_14411 = ~n_14406 &  n_14410;
assign n_14412 =  n_13869 & ~n_14411;
assign n_14413 = ~n_14409 &  n_14412;
assign n_14414 = ~n_14401 & ~n_14413;
assign n_14415 = ~n_14400 &  n_14414;
assign n_14416 =  x_792 & ~n_14415;
assign n_14417 = ~x_792 &  n_14415;
assign n_14418 = ~n_14416 & ~n_14417;
assign n_14419 = ~x_2711 &  n_14389;
assign n_14420 =  x_2711 & ~n_14389;
assign n_14421 = ~n_14419 & ~n_14420;
assign n_14422 = ~n_14393 & ~n_14397;
assign n_14423 =  n_14421 & ~n_14422;
assign n_14424 = ~n_14421 &  n_14422;
assign n_14425 = ~n_14423 & ~n_14424;
assign n_14426 = ~x_2295 & ~n_14425;
assign n_14427 =  x_2295 & ~n_14424;
assign n_14428 = ~n_14423 &  n_14427;
assign n_14429 =  n_13860 & ~n_14428;
assign n_14430 = ~n_14426 &  n_14429;
assign n_14431 =  x_791 & ~n_13866;
assign n_14432 = ~x_471 &  n_14402;
assign n_14433 =  x_471 & ~n_14402;
assign n_14434 = ~n_14432 & ~n_14433;
assign n_14435 = ~n_14406 & ~n_14410;
assign n_14436 =  n_14434 & ~n_14435;
assign n_14437 = ~n_14434 &  n_14435;
assign n_14438 = ~n_14436 & ~n_14437;
assign n_14439 = ~x_1207 & ~n_14438;
assign n_14440 =  x_1207 & ~n_14437;
assign n_14441 = ~n_14436 &  n_14440;
assign n_14442 =  n_13869 & ~n_14441;
assign n_14443 = ~n_14439 &  n_14442;
assign n_14444 = ~n_14431 & ~n_14443;
assign n_14445 = ~n_14430 &  n_14444;
assign n_14446 =  x_791 & ~n_14445;
assign n_14447 = ~x_791 &  n_14445;
assign n_14448 = ~n_14446 & ~n_14447;
assign n_14449 = ~x_2710 &  n_14419;
assign n_14450 =  x_2710 & ~n_14419;
assign n_14451 = ~n_14449 & ~n_14450;
assign n_14452 = ~n_14423 & ~n_14427;
assign n_14453 =  n_14451 & ~n_14452;
assign n_14454 = ~n_14451 &  n_14452;
assign n_14455 = ~n_14453 & ~n_14454;
assign n_14456 = ~x_2294 & ~n_14455;
assign n_14457 =  x_2294 & ~n_14454;
assign n_14458 = ~n_14453 &  n_14457;
assign n_14459 =  n_13860 & ~n_14458;
assign n_14460 = ~n_14456 &  n_14459;
assign n_14461 =  x_790 & ~n_13866;
assign n_14462 = ~x_470 &  n_14432;
assign n_14463 =  x_470 & ~n_14432;
assign n_14464 = ~n_14462 & ~n_14463;
assign n_14465 = ~n_14436 & ~n_14440;
assign n_14466 =  n_14464 & ~n_14465;
assign n_14467 = ~n_14464 &  n_14465;
assign n_14468 = ~n_14466 & ~n_14467;
assign n_14469 = ~x_1206 & ~n_14468;
assign n_14470 =  x_1206 & ~n_14467;
assign n_14471 = ~n_14466 &  n_14470;
assign n_14472 =  n_13869 & ~n_14471;
assign n_14473 = ~n_14469 &  n_14472;
assign n_14474 = ~n_14461 & ~n_14473;
assign n_14475 = ~n_14460 &  n_14474;
assign n_14476 =  x_790 & ~n_14475;
assign n_14477 = ~x_790 &  n_14475;
assign n_14478 = ~n_14476 & ~n_14477;
assign n_14479 = ~x_2709 &  n_14449;
assign n_14480 =  x_2709 & ~n_14449;
assign n_14481 = ~n_14479 & ~n_14480;
assign n_14482 = ~n_14453 & ~n_14457;
assign n_14483 =  n_14481 & ~n_14482;
assign n_14484 = ~n_14481 &  n_14482;
assign n_14485 = ~n_14483 & ~n_14484;
assign n_14486 = ~x_2293 & ~n_14485;
assign n_14487 =  x_2293 & ~n_14484;
assign n_14488 = ~n_14483 &  n_14487;
assign n_14489 =  n_13860 & ~n_14488;
assign n_14490 = ~n_14486 &  n_14489;
assign n_14491 =  x_789 & ~n_13866;
assign n_14492 = ~x_469 &  n_14462;
assign n_14493 =  x_469 & ~n_14462;
assign n_14494 = ~n_14492 & ~n_14493;
assign n_14495 = ~n_14466 & ~n_14470;
assign n_14496 =  n_14494 & ~n_14495;
assign n_14497 = ~n_14494 &  n_14495;
assign n_14498 = ~n_14496 & ~n_14497;
assign n_14499 = ~x_1205 & ~n_14498;
assign n_14500 =  x_1205 & ~n_14497;
assign n_14501 = ~n_14496 &  n_14500;
assign n_14502 =  n_13869 & ~n_14501;
assign n_14503 = ~n_14499 &  n_14502;
assign n_14504 = ~n_14491 & ~n_14503;
assign n_14505 = ~n_14490 &  n_14504;
assign n_14506 =  x_789 & ~n_14505;
assign n_14507 = ~x_789 &  n_14505;
assign n_14508 = ~n_14506 & ~n_14507;
assign n_14509 = ~x_2708 &  n_14479;
assign n_14510 =  x_2708 & ~n_14479;
assign n_14511 = ~n_14509 & ~n_14510;
assign n_14512 = ~n_14483 & ~n_14487;
assign n_14513 =  n_14511 & ~n_14512;
assign n_14514 = ~n_14511 &  n_14512;
assign n_14515 = ~n_14513 & ~n_14514;
assign n_14516 = ~x_2292 & ~n_14515;
assign n_14517 =  x_2292 & ~n_14514;
assign n_14518 = ~n_14513 &  n_14517;
assign n_14519 =  n_13860 & ~n_14518;
assign n_14520 = ~n_14516 &  n_14519;
assign n_14521 =  x_788 & ~n_13866;
assign n_14522 = ~x_468 &  n_14492;
assign n_14523 =  x_468 & ~n_14492;
assign n_14524 = ~n_14522 & ~n_14523;
assign n_14525 = ~n_14496 & ~n_14500;
assign n_14526 =  n_14524 & ~n_14525;
assign n_14527 = ~n_14524 &  n_14525;
assign n_14528 = ~n_14526 & ~n_14527;
assign n_14529 = ~x_1204 & ~n_14528;
assign n_14530 =  x_1204 & ~n_14527;
assign n_14531 = ~n_14526 &  n_14530;
assign n_14532 =  n_13869 & ~n_14531;
assign n_14533 = ~n_14529 &  n_14532;
assign n_14534 = ~n_14521 & ~n_14533;
assign n_14535 = ~n_14520 &  n_14534;
assign n_14536 =  x_788 & ~n_14535;
assign n_14537 = ~x_788 &  n_14535;
assign n_14538 = ~n_14536 & ~n_14537;
assign n_14539 = ~x_2707 &  n_14509;
assign n_14540 =  x_2707 & ~n_14509;
assign n_14541 = ~n_14539 & ~n_14540;
assign n_14542 = ~n_14513 & ~n_14517;
assign n_14543 =  n_14541 & ~n_14542;
assign n_14544 = ~n_14541 &  n_14542;
assign n_14545 = ~n_14543 & ~n_14544;
assign n_14546 = ~x_2291 & ~n_14545;
assign n_14547 =  x_2291 & ~n_14544;
assign n_14548 = ~n_14543 &  n_14547;
assign n_14549 =  n_13860 & ~n_14548;
assign n_14550 = ~n_14546 &  n_14549;
assign n_14551 =  x_787 & ~n_13866;
assign n_14552 = ~x_467 &  n_14522;
assign n_14553 =  x_467 & ~n_14522;
assign n_14554 = ~n_14552 & ~n_14553;
assign n_14555 = ~n_14526 & ~n_14530;
assign n_14556 =  n_14554 & ~n_14555;
assign n_14557 = ~n_14554 &  n_14555;
assign n_14558 = ~n_14556 & ~n_14557;
assign n_14559 = ~x_1203 & ~n_14558;
assign n_14560 =  x_1203 & ~n_14557;
assign n_14561 = ~n_14556 &  n_14560;
assign n_14562 =  n_13869 & ~n_14561;
assign n_14563 = ~n_14559 &  n_14562;
assign n_14564 = ~n_14551 & ~n_14563;
assign n_14565 = ~n_14550 &  n_14564;
assign n_14566 =  x_787 & ~n_14565;
assign n_14567 = ~x_787 &  n_14565;
assign n_14568 = ~n_14566 & ~n_14567;
assign n_14569 = ~x_2706 &  n_14539;
assign n_14570 =  x_2706 & ~n_14539;
assign n_14571 = ~n_14569 & ~n_14570;
assign n_14572 = ~n_14543 & ~n_14547;
assign n_14573 =  n_14571 & ~n_14572;
assign n_14574 = ~n_14571 &  n_14572;
assign n_14575 = ~n_14573 & ~n_14574;
assign n_14576 = ~x_2290 & ~n_14575;
assign n_14577 =  x_2290 & ~n_14574;
assign n_14578 = ~n_14573 &  n_14577;
assign n_14579 =  n_13860 & ~n_14578;
assign n_14580 = ~n_14576 &  n_14579;
assign n_14581 =  x_786 & ~n_13866;
assign n_14582 = ~x_466 &  n_14552;
assign n_14583 =  x_466 & ~n_14552;
assign n_14584 = ~n_14582 & ~n_14583;
assign n_14585 = ~n_14556 & ~n_14560;
assign n_14586 =  n_14584 & ~n_14585;
assign n_14587 = ~n_14584 &  n_14585;
assign n_14588 = ~n_14586 & ~n_14587;
assign n_14589 = ~x_1202 & ~n_14588;
assign n_14590 =  x_1202 & ~n_14587;
assign n_14591 = ~n_14586 &  n_14590;
assign n_14592 =  n_13869 & ~n_14591;
assign n_14593 = ~n_14589 &  n_14592;
assign n_14594 = ~n_14581 & ~n_14593;
assign n_14595 = ~n_14580 &  n_14594;
assign n_14596 =  x_786 & ~n_14595;
assign n_14597 = ~x_786 &  n_14595;
assign n_14598 = ~n_14596 & ~n_14597;
assign n_14599 = ~x_2705 &  n_14569;
assign n_14600 =  x_2705 & ~n_14569;
assign n_14601 = ~n_14599 & ~n_14600;
assign n_14602 = ~n_14573 & ~n_14577;
assign n_14603 =  n_14601 & ~n_14602;
assign n_14604 = ~n_14601 &  n_14602;
assign n_14605 = ~n_14603 & ~n_14604;
assign n_14606 = ~x_2289 & ~n_14605;
assign n_14607 =  x_2289 & ~n_14604;
assign n_14608 = ~n_14603 &  n_14607;
assign n_14609 =  n_13860 & ~n_14608;
assign n_14610 = ~n_14606 &  n_14609;
assign n_14611 =  x_785 & ~n_13866;
assign n_14612 = ~x_465 &  n_14582;
assign n_14613 =  x_465 & ~n_14582;
assign n_14614 = ~n_14612 & ~n_14613;
assign n_14615 = ~n_14586 & ~n_14590;
assign n_14616 =  n_14614 & ~n_14615;
assign n_14617 = ~n_14614 &  n_14615;
assign n_14618 = ~n_14616 & ~n_14617;
assign n_14619 = ~x_1201 & ~n_14618;
assign n_14620 =  x_1201 & ~n_14617;
assign n_14621 = ~n_14616 &  n_14620;
assign n_14622 =  n_13869 & ~n_14621;
assign n_14623 = ~n_14619 &  n_14622;
assign n_14624 = ~n_14611 & ~n_14623;
assign n_14625 = ~n_14610 &  n_14624;
assign n_14626 =  x_785 & ~n_14625;
assign n_14627 = ~x_785 &  n_14625;
assign n_14628 = ~n_14626 & ~n_14627;
assign n_14629 = ~x_2704 &  n_14599;
assign n_14630 =  x_2704 & ~n_14599;
assign n_14631 = ~n_14629 & ~n_14630;
assign n_14632 = ~n_14603 & ~n_14607;
assign n_14633 =  n_14631 & ~n_14632;
assign n_14634 = ~n_14631 &  n_14632;
assign n_14635 = ~n_14633 & ~n_14634;
assign n_14636 = ~x_2288 & ~n_14635;
assign n_14637 =  x_2288 & ~n_14634;
assign n_14638 = ~n_14633 &  n_14637;
assign n_14639 =  n_13860 & ~n_14638;
assign n_14640 = ~n_14636 &  n_14639;
assign n_14641 =  x_784 & ~n_13866;
assign n_14642 = ~x_464 &  n_14612;
assign n_14643 =  x_464 & ~n_14612;
assign n_14644 = ~n_14642 & ~n_14643;
assign n_14645 = ~n_14616 & ~n_14620;
assign n_14646 =  n_14644 & ~n_14645;
assign n_14647 = ~n_14644 &  n_14645;
assign n_14648 = ~n_14646 & ~n_14647;
assign n_14649 = ~x_1200 & ~n_14648;
assign n_14650 =  x_1200 & ~n_14647;
assign n_14651 = ~n_14646 &  n_14650;
assign n_14652 =  n_13869 & ~n_14651;
assign n_14653 = ~n_14649 &  n_14652;
assign n_14654 = ~n_14641 & ~n_14653;
assign n_14655 = ~n_14640 &  n_14654;
assign n_14656 =  x_784 & ~n_14655;
assign n_14657 = ~x_784 &  n_14655;
assign n_14658 = ~n_14656 & ~n_14657;
assign n_14659 = ~x_2703 &  n_14629;
assign n_14660 =  x_2703 & ~n_14629;
assign n_14661 = ~n_14659 & ~n_14660;
assign n_14662 = ~n_14633 & ~n_14637;
assign n_14663 =  n_14661 & ~n_14662;
assign n_14664 = ~n_14661 &  n_14662;
assign n_14665 = ~n_14663 & ~n_14664;
assign n_14666 = ~x_2287 & ~n_14665;
assign n_14667 =  x_2287 & ~n_14664;
assign n_14668 = ~n_14663 &  n_14667;
assign n_14669 =  n_13860 & ~n_14668;
assign n_14670 = ~n_14666 &  n_14669;
assign n_14671 =  x_783 & ~n_13866;
assign n_14672 = ~x_463 &  n_14642;
assign n_14673 =  x_463 & ~n_14642;
assign n_14674 = ~n_14672 & ~n_14673;
assign n_14675 = ~n_14646 & ~n_14650;
assign n_14676 =  n_14674 & ~n_14675;
assign n_14677 = ~n_14674 &  n_14675;
assign n_14678 = ~n_14676 & ~n_14677;
assign n_14679 = ~x_1199 & ~n_14678;
assign n_14680 =  x_1199 & ~n_14677;
assign n_14681 = ~n_14676 &  n_14680;
assign n_14682 =  n_13869 & ~n_14681;
assign n_14683 = ~n_14679 &  n_14682;
assign n_14684 = ~n_14671 & ~n_14683;
assign n_14685 = ~n_14670 &  n_14684;
assign n_14686 =  x_783 & ~n_14685;
assign n_14687 = ~x_783 &  n_14685;
assign n_14688 = ~n_14686 & ~n_14687;
assign n_14689 = ~x_2702 &  n_14659;
assign n_14690 =  x_2702 & ~n_14659;
assign n_14691 = ~n_14689 & ~n_14690;
assign n_14692 = ~n_14663 & ~n_14667;
assign n_14693 =  n_14691 & ~n_14692;
assign n_14694 = ~n_14691 &  n_14692;
assign n_14695 = ~n_14693 & ~n_14694;
assign n_14696 = ~x_2286 & ~n_14695;
assign n_14697 =  x_2286 & ~n_14694;
assign n_14698 = ~n_14693 &  n_14697;
assign n_14699 =  n_13860 & ~n_14698;
assign n_14700 = ~n_14696 &  n_14699;
assign n_14701 =  x_782 & ~n_13866;
assign n_14702 = ~x_462 &  n_14672;
assign n_14703 =  x_462 & ~n_14672;
assign n_14704 = ~n_14702 & ~n_14703;
assign n_14705 = ~n_14676 & ~n_14680;
assign n_14706 =  n_14704 & ~n_14705;
assign n_14707 = ~n_14704 &  n_14705;
assign n_14708 = ~n_14706 & ~n_14707;
assign n_14709 = ~x_1198 & ~n_14708;
assign n_14710 =  x_1198 & ~n_14707;
assign n_14711 = ~n_14706 &  n_14710;
assign n_14712 =  n_13869 & ~n_14711;
assign n_14713 = ~n_14709 &  n_14712;
assign n_14714 = ~n_14701 & ~n_14713;
assign n_14715 = ~n_14700 &  n_14714;
assign n_14716 =  x_782 & ~n_14715;
assign n_14717 = ~x_782 &  n_14715;
assign n_14718 = ~n_14716 & ~n_14717;
assign n_14719 = ~x_2701 &  n_14689;
assign n_14720 =  x_2701 & ~n_14689;
assign n_14721 = ~n_14719 & ~n_14720;
assign n_14722 = ~n_14693 & ~n_14697;
assign n_14723 =  n_14721 & ~n_14722;
assign n_14724 = ~n_14721 &  n_14722;
assign n_14725 = ~n_14723 & ~n_14724;
assign n_14726 = ~x_2285 & ~n_14725;
assign n_14727 =  x_2285 & ~n_14724;
assign n_14728 = ~n_14723 &  n_14727;
assign n_14729 =  n_13860 & ~n_14728;
assign n_14730 = ~n_14726 &  n_14729;
assign n_14731 =  x_781 & ~n_13866;
assign n_14732 = ~x_461 &  n_14702;
assign n_14733 =  x_461 & ~n_14702;
assign n_14734 = ~n_14732 & ~n_14733;
assign n_14735 = ~n_14706 & ~n_14710;
assign n_14736 =  n_14734 & ~n_14735;
assign n_14737 = ~n_14734 &  n_14735;
assign n_14738 = ~n_14736 & ~n_14737;
assign n_14739 = ~x_1197 & ~n_14738;
assign n_14740 =  x_1197 & ~n_14737;
assign n_14741 = ~n_14736 &  n_14740;
assign n_14742 =  n_13869 & ~n_14741;
assign n_14743 = ~n_14739 &  n_14742;
assign n_14744 = ~n_14731 & ~n_14743;
assign n_14745 = ~n_14730 &  n_14744;
assign n_14746 =  x_781 & ~n_14745;
assign n_14747 = ~x_781 &  n_14745;
assign n_14748 = ~n_14746 & ~n_14747;
assign n_14749 = ~x_2700 &  n_14719;
assign n_14750 =  x_2700 & ~n_14719;
assign n_14751 = ~n_14749 & ~n_14750;
assign n_14752 = ~n_14723 & ~n_14727;
assign n_14753 =  n_14751 & ~n_14752;
assign n_14754 = ~n_14751 &  n_14752;
assign n_14755 = ~n_14753 & ~n_14754;
assign n_14756 = ~x_2284 & ~n_14755;
assign n_14757 =  x_2284 & ~n_14754;
assign n_14758 = ~n_14753 &  n_14757;
assign n_14759 =  n_13860 & ~n_14758;
assign n_14760 = ~n_14756 &  n_14759;
assign n_14761 =  x_780 & ~n_13866;
assign n_14762 = ~x_460 &  n_14732;
assign n_14763 =  x_460 & ~n_14732;
assign n_14764 = ~n_14762 & ~n_14763;
assign n_14765 = ~n_14736 & ~n_14740;
assign n_14766 =  n_14764 & ~n_14765;
assign n_14767 = ~n_14764 &  n_14765;
assign n_14768 = ~n_14766 & ~n_14767;
assign n_14769 = ~x_1196 & ~n_14768;
assign n_14770 =  x_1196 & ~n_14767;
assign n_14771 = ~n_14766 &  n_14770;
assign n_14772 =  n_13869 & ~n_14771;
assign n_14773 = ~n_14769 &  n_14772;
assign n_14774 = ~n_14761 & ~n_14773;
assign n_14775 = ~n_14760 &  n_14774;
assign n_14776 =  x_780 & ~n_14775;
assign n_14777 = ~x_780 &  n_14775;
assign n_14778 = ~n_14776 & ~n_14777;
assign n_14779 = ~n_14766 & ~n_14770;
assign n_14780 =  x_459 & ~x_1195;
assign n_14781 = ~x_459 &  x_1195;
assign n_14782 = ~n_14780 & ~n_14781;
assign n_14783 =  n_14762 &  n_14782;
assign n_14784 = ~n_14762 & ~n_14782;
assign n_14785 = ~n_14783 & ~n_14784;
assign n_14786 =  n_14779 & ~n_14785;
assign n_14787 = ~n_14779 &  n_14785;
assign n_14788 =  n_13869 & ~n_14787;
assign n_14789 = ~n_14786 &  n_14788;
assign n_14790 =  x_779 & ~n_13866;
assign n_14791 = ~n_14753 & ~n_14757;
assign n_14792 =  x_2283 & ~x_2699;
assign n_14793 = ~x_2283 &  x_2699;
assign n_14794 = ~n_14792 & ~n_14793;
assign n_14795 =  n_14749 &  n_14794;
assign n_14796 = ~n_14749 & ~n_14794;
assign n_14797 = ~n_14795 & ~n_14796;
assign n_14798 =  n_14791 & ~n_14797;
assign n_14799 = ~n_14791 &  n_14797;
assign n_14800 =  n_13860 & ~n_14799;
assign n_14801 = ~n_14798 &  n_14800;
assign n_14802 = ~n_14790 & ~n_14801;
assign n_14803 = ~n_14789 &  n_14802;
assign n_14804 =  x_779 & ~n_14803;
assign n_14805 = ~x_779 &  n_14803;
assign n_14806 = ~n_14804 & ~n_14805;
assign n_14807 =  n_2100 &  n_7;
assign n_14808 =  x_39 &  n_14807;
assign n_14809 = ~n_8 & ~n_14808;
assign n_14810 =  n_586 & ~n_14809;
assign n_14811 =  x_778 & ~n_14810;
assign n_14812 =  n_8818 &  n_8;
assign n_14813 =  x_714 &  x_1930;
assign n_14814 = ~x_714 & ~x_1930;
assign n_14815 = ~n_14813 & ~n_14814;
assign n_14816 =  n_14812 &  n_14815;
assign n_14817 =  n_8 &  n_587;
assign n_14818 =  x_2378 &  x_2666;
assign n_14819 = ~x_2378 & ~x_2666;
assign n_14820 = ~n_14818 & ~n_14819;
assign n_14821 =  n_14817 &  n_14820;
assign n_14822 = ~n_14816 & ~n_14821;
assign n_14823 = ~n_14811 &  n_14822;
assign n_14824 =  x_778 & ~n_14823;
assign n_14825 = ~x_778 &  n_14823;
assign n_14826 = ~n_14824 & ~n_14825;
assign n_14827 =  x_777 & ~n_14810;
assign n_14828 = ~x_1929 & ~x_1930;
assign n_14829 =  x_1929 &  x_1930;
assign n_14830 = ~n_14828 & ~n_14829;
assign n_14831 =  x_713 &  n_14830;
assign n_14832 = ~x_713 & ~n_14830;
assign n_14833 = ~n_14831 & ~n_14832;
assign n_14834 = ~n_14813 & ~n_14833;
assign n_14835 =  n_14813 &  n_14833;
assign n_14836 =  n_14812 & ~n_14835;
assign n_14837 = ~n_14834 &  n_14836;
assign n_14838 = ~x_2665 & ~x_2666;
assign n_14839 =  x_2665 &  x_2666;
assign n_14840 = ~n_14838 & ~n_14839;
assign n_14841 =  x_2377 &  n_14840;
assign n_14842 = ~x_2377 & ~n_14840;
assign n_14843 = ~n_14841 & ~n_14842;
assign n_14844 = ~n_14818 & ~n_14843;
assign n_14845 =  n_14818 &  n_14843;
assign n_14846 =  n_14817 & ~n_14845;
assign n_14847 = ~n_14844 &  n_14846;
assign n_14848 = ~n_14837 & ~n_14847;
assign n_14849 = ~n_14827 &  n_14848;
assign n_14850 =  x_777 & ~n_14849;
assign n_14851 = ~x_777 &  n_14849;
assign n_14852 = ~n_14850 & ~n_14851;
assign n_14853 = ~x_1928 &  n_14828;
assign n_14854 =  x_1928 & ~n_14828;
assign n_14855 = ~n_14853 & ~n_14854;
assign n_14856 = ~x_713 &  x_1929;
assign n_14857 =  n_14813 & ~n_14856;
assign n_14858 = ~n_14857 & ~n_14831;
assign n_14859 =  n_14855 & ~n_14858;
assign n_14860 = ~n_14855 &  n_14858;
assign n_14861 = ~n_14859 & ~n_14860;
assign n_14862 = ~x_712 & ~n_14861;
assign n_14863 =  x_712 & ~n_14860;
assign n_14864 = ~n_14859 &  n_14863;
assign n_14865 =  n_14812 & ~n_14864;
assign n_14866 = ~n_14862 &  n_14865;
assign n_14867 =  x_776 & ~n_14810;
assign n_14868 = ~x_2664 &  n_14838;
assign n_14869 =  x_2664 & ~n_14838;
assign n_14870 = ~n_14868 & ~n_14869;
assign n_14871 = ~x_2377 &  x_2665;
assign n_14872 =  n_14818 & ~n_14871;
assign n_14873 = ~n_14872 & ~n_14841;
assign n_14874 =  n_14870 & ~n_14873;
assign n_14875 = ~n_14870 &  n_14873;
assign n_14876 = ~n_14874 & ~n_14875;
assign n_14877 = ~x_2376 & ~n_14876;
assign n_14878 =  x_2376 & ~n_14875;
assign n_14879 = ~n_14874 &  n_14878;
assign n_14880 =  n_14817 & ~n_14879;
assign n_14881 = ~n_14877 &  n_14880;
assign n_14882 = ~n_14867 & ~n_14881;
assign n_14883 = ~n_14866 &  n_14882;
assign n_14884 =  x_776 & ~n_14883;
assign n_14885 = ~x_776 &  n_14883;
assign n_14886 = ~n_14884 & ~n_14885;
assign n_14887 = ~x_2663 &  n_14868;
assign n_14888 =  x_2663 & ~n_14868;
assign n_14889 = ~n_14887 & ~n_14888;
assign n_14890 = ~n_14874 & ~n_14878;
assign n_14891 =  n_14889 & ~n_14890;
assign n_14892 = ~n_14889 &  n_14890;
assign n_14893 = ~n_14891 & ~n_14892;
assign n_14894 = ~x_2375 & ~n_14893;
assign n_14895 =  x_2375 & ~n_14892;
assign n_14896 = ~n_14891 &  n_14895;
assign n_14897 =  n_14817 & ~n_14896;
assign n_14898 = ~n_14894 &  n_14897;
assign n_14899 =  x_775 & ~n_14810;
assign n_14900 = ~x_1927 &  n_14853;
assign n_14901 =  x_1927 & ~n_14853;
assign n_14902 = ~n_14900 & ~n_14901;
assign n_14903 = ~n_14859 & ~n_14863;
assign n_14904 =  n_14902 & ~n_14903;
assign n_14905 = ~n_14902 &  n_14903;
assign n_14906 = ~n_14904 & ~n_14905;
assign n_14907 = ~x_711 & ~n_14906;
assign n_14908 =  x_711 & ~n_14905;
assign n_14909 = ~n_14904 &  n_14908;
assign n_14910 =  n_14812 & ~n_14909;
assign n_14911 = ~n_14907 &  n_14910;
assign n_14912 = ~n_14899 & ~n_14911;
assign n_14913 = ~n_14898 &  n_14912;
assign n_14914 =  x_775 & ~n_14913;
assign n_14915 = ~x_775 &  n_14913;
assign n_14916 = ~n_14914 & ~n_14915;
assign n_14917 = ~x_2662 &  n_14887;
assign n_14918 =  x_2662 & ~n_14887;
assign n_14919 = ~n_14917 & ~n_14918;
assign n_14920 = ~n_14891 & ~n_14895;
assign n_14921 =  n_14919 & ~n_14920;
assign n_14922 = ~n_14919 &  n_14920;
assign n_14923 = ~n_14921 & ~n_14922;
assign n_14924 = ~x_2374 & ~n_14923;
assign n_14925 =  x_2374 & ~n_14922;
assign n_14926 = ~n_14921 &  n_14925;
assign n_14927 =  n_14817 & ~n_14926;
assign n_14928 = ~n_14924 &  n_14927;
assign n_14929 =  x_774 & ~n_14810;
assign n_14930 = ~x_1926 &  n_14900;
assign n_14931 =  x_1926 & ~n_14900;
assign n_14932 = ~n_14930 & ~n_14931;
assign n_14933 = ~n_14904 & ~n_14908;
assign n_14934 =  n_14932 & ~n_14933;
assign n_14935 = ~n_14932 &  n_14933;
assign n_14936 = ~n_14934 & ~n_14935;
assign n_14937 = ~x_710 & ~n_14936;
assign n_14938 =  x_710 & ~n_14935;
assign n_14939 = ~n_14934 &  n_14938;
assign n_14940 =  n_14812 & ~n_14939;
assign n_14941 = ~n_14937 &  n_14940;
assign n_14942 = ~n_14929 & ~n_14941;
assign n_14943 = ~n_14928 &  n_14942;
assign n_14944 =  x_774 & ~n_14943;
assign n_14945 = ~x_774 &  n_14943;
assign n_14946 = ~n_14944 & ~n_14945;
assign n_14947 = ~x_2661 &  n_14917;
assign n_14948 =  x_2661 & ~n_14917;
assign n_14949 = ~n_14947 & ~n_14948;
assign n_14950 = ~n_14921 & ~n_14925;
assign n_14951 =  n_14949 & ~n_14950;
assign n_14952 = ~n_14949 &  n_14950;
assign n_14953 = ~n_14951 & ~n_14952;
assign n_14954 = ~x_2373 & ~n_14953;
assign n_14955 =  x_2373 & ~n_14952;
assign n_14956 = ~n_14951 &  n_14955;
assign n_14957 =  n_14817 & ~n_14956;
assign n_14958 = ~n_14954 &  n_14957;
assign n_14959 =  x_773 & ~n_14810;
assign n_14960 = ~x_1925 &  n_14930;
assign n_14961 =  x_1925 & ~n_14930;
assign n_14962 = ~n_14960 & ~n_14961;
assign n_14963 = ~n_14934 & ~n_14938;
assign n_14964 =  n_14962 & ~n_14963;
assign n_14965 = ~n_14962 &  n_14963;
assign n_14966 = ~n_14964 & ~n_14965;
assign n_14967 = ~x_709 & ~n_14966;
assign n_14968 =  x_709 & ~n_14965;
assign n_14969 = ~n_14964 &  n_14968;
assign n_14970 =  n_14812 & ~n_14969;
assign n_14971 = ~n_14967 &  n_14970;
assign n_14972 = ~n_14959 & ~n_14971;
assign n_14973 = ~n_14958 &  n_14972;
assign n_14974 =  x_773 & ~n_14973;
assign n_14975 = ~x_773 &  n_14973;
assign n_14976 = ~n_14974 & ~n_14975;
assign n_14977 = ~x_2660 &  n_14947;
assign n_14978 =  x_2660 & ~n_14947;
assign n_14979 = ~n_14977 & ~n_14978;
assign n_14980 = ~n_14951 & ~n_14955;
assign n_14981 =  n_14979 & ~n_14980;
assign n_14982 = ~n_14979 &  n_14980;
assign n_14983 = ~n_14981 & ~n_14982;
assign n_14984 = ~x_2372 & ~n_14983;
assign n_14985 =  x_2372 & ~n_14982;
assign n_14986 = ~n_14981 &  n_14985;
assign n_14987 =  n_14817 & ~n_14986;
assign n_14988 = ~n_14984 &  n_14987;
assign n_14989 =  x_772 & ~n_14810;
assign n_14990 = ~x_1924 &  n_14960;
assign n_14991 =  x_1924 & ~n_14960;
assign n_14992 = ~n_14990 & ~n_14991;
assign n_14993 = ~n_14964 & ~n_14968;
assign n_14994 =  n_14992 & ~n_14993;
assign n_14995 = ~n_14992 &  n_14993;
assign n_14996 = ~n_14994 & ~n_14995;
assign n_14997 = ~x_708 & ~n_14996;
assign n_14998 =  x_708 & ~n_14995;
assign n_14999 = ~n_14994 &  n_14998;
assign n_15000 =  n_14812 & ~n_14999;
assign n_15001 = ~n_14997 &  n_15000;
assign n_15002 = ~n_14989 & ~n_15001;
assign n_15003 = ~n_14988 &  n_15002;
assign n_15004 =  x_772 & ~n_15003;
assign n_15005 = ~x_772 &  n_15003;
assign n_15006 = ~n_15004 & ~n_15005;
assign n_15007 = ~x_2659 &  n_14977;
assign n_15008 =  x_2659 & ~n_14977;
assign n_15009 = ~n_15007 & ~n_15008;
assign n_15010 = ~n_14981 & ~n_14985;
assign n_15011 =  n_15009 & ~n_15010;
assign n_15012 = ~n_15009 &  n_15010;
assign n_15013 = ~n_15011 & ~n_15012;
assign n_15014 = ~x_2371 & ~n_15013;
assign n_15015 =  x_2371 & ~n_15012;
assign n_15016 = ~n_15011 &  n_15015;
assign n_15017 =  n_14817 & ~n_15016;
assign n_15018 = ~n_15014 &  n_15017;
assign n_15019 =  x_771 & ~n_14810;
assign n_15020 = ~x_1923 &  n_14990;
assign n_15021 =  x_1923 & ~n_14990;
assign n_15022 = ~n_15020 & ~n_15021;
assign n_15023 = ~n_14994 & ~n_14998;
assign n_15024 =  n_15022 & ~n_15023;
assign n_15025 = ~n_15022 &  n_15023;
assign n_15026 = ~n_15024 & ~n_15025;
assign n_15027 = ~x_707 & ~n_15026;
assign n_15028 =  x_707 & ~n_15025;
assign n_15029 = ~n_15024 &  n_15028;
assign n_15030 =  n_14812 & ~n_15029;
assign n_15031 = ~n_15027 &  n_15030;
assign n_15032 = ~n_15019 & ~n_15031;
assign n_15033 = ~n_15018 &  n_15032;
assign n_15034 =  x_771 & ~n_15033;
assign n_15035 = ~x_771 &  n_15033;
assign n_15036 = ~n_15034 & ~n_15035;
assign n_15037 = ~x_2658 &  n_15007;
assign n_15038 =  x_2658 & ~n_15007;
assign n_15039 = ~n_15037 & ~n_15038;
assign n_15040 = ~n_15011 & ~n_15015;
assign n_15041 =  n_15039 & ~n_15040;
assign n_15042 = ~n_15039 &  n_15040;
assign n_15043 = ~n_15041 & ~n_15042;
assign n_15044 = ~x_2370 & ~n_15043;
assign n_15045 =  x_2370 & ~n_15042;
assign n_15046 = ~n_15041 &  n_15045;
assign n_15047 =  n_14817 & ~n_15046;
assign n_15048 = ~n_15044 &  n_15047;
assign n_15049 =  x_770 & ~n_14810;
assign n_15050 = ~x_1922 &  n_15020;
assign n_15051 =  x_1922 & ~n_15020;
assign n_15052 = ~n_15050 & ~n_15051;
assign n_15053 = ~n_15024 & ~n_15028;
assign n_15054 =  n_15052 & ~n_15053;
assign n_15055 = ~n_15052 &  n_15053;
assign n_15056 = ~n_15054 & ~n_15055;
assign n_15057 = ~x_706 & ~n_15056;
assign n_15058 =  x_706 & ~n_15055;
assign n_15059 = ~n_15054 &  n_15058;
assign n_15060 =  n_14812 & ~n_15059;
assign n_15061 = ~n_15057 &  n_15060;
assign n_15062 = ~n_15049 & ~n_15061;
assign n_15063 = ~n_15048 &  n_15062;
assign n_15064 =  x_770 & ~n_15063;
assign n_15065 = ~x_770 &  n_15063;
assign n_15066 = ~n_15064 & ~n_15065;
assign n_15067 = ~x_2657 &  n_15037;
assign n_15068 =  x_2657 & ~n_15037;
assign n_15069 = ~n_15067 & ~n_15068;
assign n_15070 = ~n_15041 & ~n_15045;
assign n_15071 =  n_15069 & ~n_15070;
assign n_15072 = ~n_15069 &  n_15070;
assign n_15073 = ~n_15071 & ~n_15072;
assign n_15074 = ~x_2369 & ~n_15073;
assign n_15075 =  x_2369 & ~n_15072;
assign n_15076 = ~n_15071 &  n_15075;
assign n_15077 =  n_14817 & ~n_15076;
assign n_15078 = ~n_15074 &  n_15077;
assign n_15079 =  x_769 & ~n_14810;
assign n_15080 = ~x_1921 &  n_15050;
assign n_15081 =  x_1921 & ~n_15050;
assign n_15082 = ~n_15080 & ~n_15081;
assign n_15083 = ~n_15054 & ~n_15058;
assign n_15084 =  n_15082 & ~n_15083;
assign n_15085 = ~n_15082 &  n_15083;
assign n_15086 = ~n_15084 & ~n_15085;
assign n_15087 = ~x_705 & ~n_15086;
assign n_15088 =  x_705 & ~n_15085;
assign n_15089 = ~n_15084 &  n_15088;
assign n_15090 =  n_14812 & ~n_15089;
assign n_15091 = ~n_15087 &  n_15090;
assign n_15092 = ~n_15079 & ~n_15091;
assign n_15093 = ~n_15078 &  n_15092;
assign n_15094 =  x_769 & ~n_15093;
assign n_15095 = ~x_769 &  n_15093;
assign n_15096 = ~n_15094 & ~n_15095;
assign n_15097 = ~x_2656 &  n_15067;
assign n_15098 =  x_2656 & ~n_15067;
assign n_15099 = ~n_15097 & ~n_15098;
assign n_15100 = ~n_15071 & ~n_15075;
assign n_15101 =  n_15099 & ~n_15100;
assign n_15102 = ~n_15099 &  n_15100;
assign n_15103 = ~n_15101 & ~n_15102;
assign n_15104 = ~x_2368 & ~n_15103;
assign n_15105 =  x_2368 & ~n_15102;
assign n_15106 = ~n_15101 &  n_15105;
assign n_15107 =  n_14817 & ~n_15106;
assign n_15108 = ~n_15104 &  n_15107;
assign n_15109 =  x_768 & ~n_14810;
assign n_15110 = ~x_1920 &  n_15080;
assign n_15111 =  x_1920 & ~n_15080;
assign n_15112 = ~n_15110 & ~n_15111;
assign n_15113 = ~n_15084 & ~n_15088;
assign n_15114 =  n_15112 & ~n_15113;
assign n_15115 = ~n_15112 &  n_15113;
assign n_15116 = ~n_15114 & ~n_15115;
assign n_15117 = ~x_704 & ~n_15116;
assign n_15118 =  x_704 & ~n_15115;
assign n_15119 = ~n_15114 &  n_15118;
assign n_15120 =  n_14812 & ~n_15119;
assign n_15121 = ~n_15117 &  n_15120;
assign n_15122 = ~n_15109 & ~n_15121;
assign n_15123 = ~n_15108 &  n_15122;
assign n_15124 =  x_768 & ~n_15123;
assign n_15125 = ~x_768 &  n_15123;
assign n_15126 = ~n_15124 & ~n_15125;
assign n_15127 = ~x_2655 &  n_15097;
assign n_15128 =  x_2655 & ~n_15097;
assign n_15129 = ~n_15127 & ~n_15128;
assign n_15130 = ~n_15101 & ~n_15105;
assign n_15131 =  n_15129 & ~n_15130;
assign n_15132 = ~n_15129 &  n_15130;
assign n_15133 = ~n_15131 & ~n_15132;
assign n_15134 = ~x_2367 & ~n_15133;
assign n_15135 =  x_2367 & ~n_15132;
assign n_15136 = ~n_15131 &  n_15135;
assign n_15137 =  n_14817 & ~n_15136;
assign n_15138 = ~n_15134 &  n_15137;
assign n_15139 =  x_767 & ~n_14810;
assign n_15140 = ~x_1919 &  n_15110;
assign n_15141 =  x_1919 & ~n_15110;
assign n_15142 = ~n_15140 & ~n_15141;
assign n_15143 = ~n_15114 & ~n_15118;
assign n_15144 =  n_15142 & ~n_15143;
assign n_15145 = ~n_15142 &  n_15143;
assign n_15146 = ~n_15144 & ~n_15145;
assign n_15147 = ~x_703 & ~n_15146;
assign n_15148 =  x_703 & ~n_15145;
assign n_15149 = ~n_15144 &  n_15148;
assign n_15150 =  n_14812 & ~n_15149;
assign n_15151 = ~n_15147 &  n_15150;
assign n_15152 = ~n_15139 & ~n_15151;
assign n_15153 = ~n_15138 &  n_15152;
assign n_15154 =  x_767 & ~n_15153;
assign n_15155 = ~x_767 &  n_15153;
assign n_15156 = ~n_15154 & ~n_15155;
assign n_15157 = ~x_2654 &  n_15127;
assign n_15158 =  x_2654 & ~n_15127;
assign n_15159 = ~n_15157 & ~n_15158;
assign n_15160 = ~n_15131 & ~n_15135;
assign n_15161 =  n_15159 & ~n_15160;
assign n_15162 = ~n_15159 &  n_15160;
assign n_15163 = ~n_15161 & ~n_15162;
assign n_15164 = ~x_2366 & ~n_15163;
assign n_15165 =  x_2366 & ~n_15162;
assign n_15166 = ~n_15161 &  n_15165;
assign n_15167 =  n_14817 & ~n_15166;
assign n_15168 = ~n_15164 &  n_15167;
assign n_15169 =  x_766 & ~n_14810;
assign n_15170 = ~x_1918 &  n_15140;
assign n_15171 =  x_1918 & ~n_15140;
assign n_15172 = ~n_15170 & ~n_15171;
assign n_15173 = ~n_15144 & ~n_15148;
assign n_15174 =  n_15172 & ~n_15173;
assign n_15175 = ~n_15172 &  n_15173;
assign n_15176 = ~n_15174 & ~n_15175;
assign n_15177 = ~x_702 & ~n_15176;
assign n_15178 =  x_702 & ~n_15175;
assign n_15179 = ~n_15174 &  n_15178;
assign n_15180 =  n_14812 & ~n_15179;
assign n_15181 = ~n_15177 &  n_15180;
assign n_15182 = ~n_15169 & ~n_15181;
assign n_15183 = ~n_15168 &  n_15182;
assign n_15184 =  x_766 & ~n_15183;
assign n_15185 = ~x_766 &  n_15183;
assign n_15186 = ~n_15184 & ~n_15185;
assign n_15187 = ~x_2653 &  n_15157;
assign n_15188 =  x_2653 & ~n_15157;
assign n_15189 = ~n_15187 & ~n_15188;
assign n_15190 = ~n_15161 & ~n_15165;
assign n_15191 =  n_15189 & ~n_15190;
assign n_15192 = ~n_15189 &  n_15190;
assign n_15193 = ~n_15191 & ~n_15192;
assign n_15194 = ~x_2365 & ~n_15193;
assign n_15195 =  x_2365 & ~n_15192;
assign n_15196 = ~n_15191 &  n_15195;
assign n_15197 =  n_14817 & ~n_15196;
assign n_15198 = ~n_15194 &  n_15197;
assign n_15199 =  x_765 & ~n_14810;
assign n_15200 = ~x_1917 &  n_15170;
assign n_15201 =  x_1917 & ~n_15170;
assign n_15202 = ~n_15200 & ~n_15201;
assign n_15203 = ~n_15174 & ~n_15178;
assign n_15204 =  n_15202 & ~n_15203;
assign n_15205 = ~n_15202 &  n_15203;
assign n_15206 = ~n_15204 & ~n_15205;
assign n_15207 = ~x_701 & ~n_15206;
assign n_15208 =  x_701 & ~n_15205;
assign n_15209 = ~n_15204 &  n_15208;
assign n_15210 =  n_14812 & ~n_15209;
assign n_15211 = ~n_15207 &  n_15210;
assign n_15212 = ~n_15199 & ~n_15211;
assign n_15213 = ~n_15198 &  n_15212;
assign n_15214 =  x_765 & ~n_15213;
assign n_15215 = ~x_765 &  n_15213;
assign n_15216 = ~n_15214 & ~n_15215;
assign n_15217 = ~x_2652 &  n_15187;
assign n_15218 =  x_2652 & ~n_15187;
assign n_15219 = ~n_15217 & ~n_15218;
assign n_15220 = ~n_15191 & ~n_15195;
assign n_15221 =  n_15219 & ~n_15220;
assign n_15222 = ~n_15219 &  n_15220;
assign n_15223 = ~n_15221 & ~n_15222;
assign n_15224 = ~x_2364 & ~n_15223;
assign n_15225 =  x_2364 & ~n_15222;
assign n_15226 = ~n_15221 &  n_15225;
assign n_15227 =  n_14817 & ~n_15226;
assign n_15228 = ~n_15224 &  n_15227;
assign n_15229 =  x_764 & ~n_14810;
assign n_15230 = ~x_1916 &  n_15200;
assign n_15231 =  x_1916 & ~n_15200;
assign n_15232 = ~n_15230 & ~n_15231;
assign n_15233 = ~n_15204 & ~n_15208;
assign n_15234 =  n_15232 & ~n_15233;
assign n_15235 = ~n_15232 &  n_15233;
assign n_15236 = ~n_15234 & ~n_15235;
assign n_15237 = ~x_700 & ~n_15236;
assign n_15238 =  x_700 & ~n_15235;
assign n_15239 = ~n_15234 &  n_15238;
assign n_15240 =  n_14812 & ~n_15239;
assign n_15241 = ~n_15237 &  n_15240;
assign n_15242 = ~n_15229 & ~n_15241;
assign n_15243 = ~n_15228 &  n_15242;
assign n_15244 =  x_764 & ~n_15243;
assign n_15245 = ~x_764 &  n_15243;
assign n_15246 = ~n_15244 & ~n_15245;
assign n_15247 = ~x_2651 &  n_15217;
assign n_15248 =  x_2651 & ~n_15217;
assign n_15249 = ~n_15247 & ~n_15248;
assign n_15250 = ~n_15221 & ~n_15225;
assign n_15251 =  n_15249 & ~n_15250;
assign n_15252 = ~n_15249 &  n_15250;
assign n_15253 = ~n_15251 & ~n_15252;
assign n_15254 = ~x_2363 & ~n_15253;
assign n_15255 =  x_2363 & ~n_15252;
assign n_15256 = ~n_15251 &  n_15255;
assign n_15257 =  n_14817 & ~n_15256;
assign n_15258 = ~n_15254 &  n_15257;
assign n_15259 =  x_763 & ~n_14810;
assign n_15260 = ~x_1915 &  n_15230;
assign n_15261 =  x_1915 & ~n_15230;
assign n_15262 = ~n_15260 & ~n_15261;
assign n_15263 = ~n_15234 & ~n_15238;
assign n_15264 =  n_15262 & ~n_15263;
assign n_15265 = ~n_15262 &  n_15263;
assign n_15266 = ~n_15264 & ~n_15265;
assign n_15267 = ~x_699 & ~n_15266;
assign n_15268 =  x_699 & ~n_15265;
assign n_15269 = ~n_15264 &  n_15268;
assign n_15270 =  n_14812 & ~n_15269;
assign n_15271 = ~n_15267 &  n_15270;
assign n_15272 = ~n_15259 & ~n_15271;
assign n_15273 = ~n_15258 &  n_15272;
assign n_15274 =  x_763 & ~n_15273;
assign n_15275 = ~x_763 &  n_15273;
assign n_15276 = ~n_15274 & ~n_15275;
assign n_15277 = ~x_2650 &  n_15247;
assign n_15278 =  x_2650 & ~n_15247;
assign n_15279 = ~n_15277 & ~n_15278;
assign n_15280 = ~n_15251 & ~n_15255;
assign n_15281 =  n_15279 & ~n_15280;
assign n_15282 = ~n_15279 &  n_15280;
assign n_15283 = ~n_15281 & ~n_15282;
assign n_15284 = ~x_2362 & ~n_15283;
assign n_15285 =  x_2362 & ~n_15282;
assign n_15286 = ~n_15281 &  n_15285;
assign n_15287 =  n_14817 & ~n_15286;
assign n_15288 = ~n_15284 &  n_15287;
assign n_15289 =  x_762 & ~n_14810;
assign n_15290 = ~x_1914 &  n_15260;
assign n_15291 =  x_1914 & ~n_15260;
assign n_15292 = ~n_15290 & ~n_15291;
assign n_15293 = ~n_15264 & ~n_15268;
assign n_15294 =  n_15292 & ~n_15293;
assign n_15295 = ~n_15292 &  n_15293;
assign n_15296 = ~n_15294 & ~n_15295;
assign n_15297 = ~x_698 & ~n_15296;
assign n_15298 =  x_698 & ~n_15295;
assign n_15299 = ~n_15294 &  n_15298;
assign n_15300 =  n_14812 & ~n_15299;
assign n_15301 = ~n_15297 &  n_15300;
assign n_15302 = ~n_15289 & ~n_15301;
assign n_15303 = ~n_15288 &  n_15302;
assign n_15304 =  x_762 & ~n_15303;
assign n_15305 = ~x_762 &  n_15303;
assign n_15306 = ~n_15304 & ~n_15305;
assign n_15307 = ~x_2649 &  n_15277;
assign n_15308 =  x_2649 & ~n_15277;
assign n_15309 = ~n_15307 & ~n_15308;
assign n_15310 = ~n_15281 & ~n_15285;
assign n_15311 =  n_15309 & ~n_15310;
assign n_15312 = ~n_15309 &  n_15310;
assign n_15313 = ~n_15311 & ~n_15312;
assign n_15314 = ~x_2361 & ~n_15313;
assign n_15315 =  x_2361 & ~n_15312;
assign n_15316 = ~n_15311 &  n_15315;
assign n_15317 =  n_14817 & ~n_15316;
assign n_15318 = ~n_15314 &  n_15317;
assign n_15319 =  x_761 & ~n_14810;
assign n_15320 = ~x_1913 &  n_15290;
assign n_15321 =  x_1913 & ~n_15290;
assign n_15322 = ~n_15320 & ~n_15321;
assign n_15323 = ~n_15294 & ~n_15298;
assign n_15324 =  n_15322 & ~n_15323;
assign n_15325 = ~n_15322 &  n_15323;
assign n_15326 = ~n_15324 & ~n_15325;
assign n_15327 = ~x_697 & ~n_15326;
assign n_15328 =  x_697 & ~n_15325;
assign n_15329 = ~n_15324 &  n_15328;
assign n_15330 =  n_14812 & ~n_15329;
assign n_15331 = ~n_15327 &  n_15330;
assign n_15332 = ~n_15319 & ~n_15331;
assign n_15333 = ~n_15318 &  n_15332;
assign n_15334 =  x_761 & ~n_15333;
assign n_15335 = ~x_761 &  n_15333;
assign n_15336 = ~n_15334 & ~n_15335;
assign n_15337 = ~x_2648 &  n_15307;
assign n_15338 =  x_2648 & ~n_15307;
assign n_15339 = ~n_15337 & ~n_15338;
assign n_15340 = ~n_15311 & ~n_15315;
assign n_15341 =  n_15339 & ~n_15340;
assign n_15342 = ~n_15339 &  n_15340;
assign n_15343 = ~n_15341 & ~n_15342;
assign n_15344 = ~x_2360 & ~n_15343;
assign n_15345 =  x_2360 & ~n_15342;
assign n_15346 = ~n_15341 &  n_15345;
assign n_15347 =  n_14817 & ~n_15346;
assign n_15348 = ~n_15344 &  n_15347;
assign n_15349 =  x_760 & ~n_14810;
assign n_15350 = ~x_1912 &  n_15320;
assign n_15351 =  x_1912 & ~n_15320;
assign n_15352 = ~n_15350 & ~n_15351;
assign n_15353 = ~n_15324 & ~n_15328;
assign n_15354 =  n_15352 & ~n_15353;
assign n_15355 = ~n_15352 &  n_15353;
assign n_15356 = ~n_15354 & ~n_15355;
assign n_15357 = ~x_696 & ~n_15356;
assign n_15358 =  x_696 & ~n_15355;
assign n_15359 = ~n_15354 &  n_15358;
assign n_15360 =  n_14812 & ~n_15359;
assign n_15361 = ~n_15357 &  n_15360;
assign n_15362 = ~n_15349 & ~n_15361;
assign n_15363 = ~n_15348 &  n_15362;
assign n_15364 =  x_760 & ~n_15363;
assign n_15365 = ~x_760 &  n_15363;
assign n_15366 = ~n_15364 & ~n_15365;
assign n_15367 = ~x_2647 &  n_15337;
assign n_15368 =  x_2647 & ~n_15337;
assign n_15369 = ~n_15367 & ~n_15368;
assign n_15370 = ~n_15341 & ~n_15345;
assign n_15371 =  n_15369 & ~n_15370;
assign n_15372 = ~n_15369 &  n_15370;
assign n_15373 = ~n_15371 & ~n_15372;
assign n_15374 = ~x_2359 & ~n_15373;
assign n_15375 =  x_2359 & ~n_15372;
assign n_15376 = ~n_15371 &  n_15375;
assign n_15377 =  n_14817 & ~n_15376;
assign n_15378 = ~n_15374 &  n_15377;
assign n_15379 =  x_759 & ~n_14810;
assign n_15380 = ~x_1911 &  n_15350;
assign n_15381 =  x_1911 & ~n_15350;
assign n_15382 = ~n_15380 & ~n_15381;
assign n_15383 = ~n_15354 & ~n_15358;
assign n_15384 =  n_15382 & ~n_15383;
assign n_15385 = ~n_15382 &  n_15383;
assign n_15386 = ~n_15384 & ~n_15385;
assign n_15387 = ~x_695 & ~n_15386;
assign n_15388 =  x_695 & ~n_15385;
assign n_15389 = ~n_15384 &  n_15388;
assign n_15390 =  n_14812 & ~n_15389;
assign n_15391 = ~n_15387 &  n_15390;
assign n_15392 = ~n_15379 & ~n_15391;
assign n_15393 = ~n_15378 &  n_15392;
assign n_15394 =  x_759 & ~n_15393;
assign n_15395 = ~x_759 &  n_15393;
assign n_15396 = ~n_15394 & ~n_15395;
assign n_15397 = ~x_2646 &  n_15367;
assign n_15398 =  x_2646 & ~n_15367;
assign n_15399 = ~n_15397 & ~n_15398;
assign n_15400 = ~n_15371 & ~n_15375;
assign n_15401 =  n_15399 & ~n_15400;
assign n_15402 = ~n_15399 &  n_15400;
assign n_15403 = ~n_15401 & ~n_15402;
assign n_15404 = ~x_2358 & ~n_15403;
assign n_15405 =  x_2358 & ~n_15402;
assign n_15406 = ~n_15401 &  n_15405;
assign n_15407 =  n_14817 & ~n_15406;
assign n_15408 = ~n_15404 &  n_15407;
assign n_15409 =  x_758 & ~n_14810;
assign n_15410 = ~x_1910 &  n_15380;
assign n_15411 =  x_1910 & ~n_15380;
assign n_15412 = ~n_15410 & ~n_15411;
assign n_15413 = ~n_15384 & ~n_15388;
assign n_15414 =  n_15412 & ~n_15413;
assign n_15415 = ~n_15412 &  n_15413;
assign n_15416 = ~n_15414 & ~n_15415;
assign n_15417 = ~x_694 & ~n_15416;
assign n_15418 =  x_694 & ~n_15415;
assign n_15419 = ~n_15414 &  n_15418;
assign n_15420 =  n_14812 & ~n_15419;
assign n_15421 = ~n_15417 &  n_15420;
assign n_15422 = ~n_15409 & ~n_15421;
assign n_15423 = ~n_15408 &  n_15422;
assign n_15424 =  x_758 & ~n_15423;
assign n_15425 = ~x_758 &  n_15423;
assign n_15426 = ~n_15424 & ~n_15425;
assign n_15427 = ~x_2645 &  n_15397;
assign n_15428 =  x_2645 & ~n_15397;
assign n_15429 = ~n_15427 & ~n_15428;
assign n_15430 = ~n_15401 & ~n_15405;
assign n_15431 =  n_15429 & ~n_15430;
assign n_15432 = ~n_15429 &  n_15430;
assign n_15433 = ~n_15431 & ~n_15432;
assign n_15434 = ~x_2357 & ~n_15433;
assign n_15435 =  x_2357 & ~n_15432;
assign n_15436 = ~n_15431 &  n_15435;
assign n_15437 =  n_14817 & ~n_15436;
assign n_15438 = ~n_15434 &  n_15437;
assign n_15439 =  x_757 & ~n_14810;
assign n_15440 = ~x_1909 &  n_15410;
assign n_15441 =  x_1909 & ~n_15410;
assign n_15442 = ~n_15440 & ~n_15441;
assign n_15443 = ~n_15414 & ~n_15418;
assign n_15444 =  n_15442 & ~n_15443;
assign n_15445 = ~n_15442 &  n_15443;
assign n_15446 = ~n_15444 & ~n_15445;
assign n_15447 = ~x_693 & ~n_15446;
assign n_15448 =  x_693 & ~n_15445;
assign n_15449 = ~n_15444 &  n_15448;
assign n_15450 =  n_14812 & ~n_15449;
assign n_15451 = ~n_15447 &  n_15450;
assign n_15452 = ~n_15439 & ~n_15451;
assign n_15453 = ~n_15438 &  n_15452;
assign n_15454 =  x_757 & ~n_15453;
assign n_15455 = ~x_757 &  n_15453;
assign n_15456 = ~n_15454 & ~n_15455;
assign n_15457 = ~x_2644 &  n_15427;
assign n_15458 =  x_2644 & ~n_15427;
assign n_15459 = ~n_15457 & ~n_15458;
assign n_15460 = ~n_15431 & ~n_15435;
assign n_15461 =  n_15459 & ~n_15460;
assign n_15462 = ~n_15459 &  n_15460;
assign n_15463 = ~n_15461 & ~n_15462;
assign n_15464 = ~x_2356 & ~n_15463;
assign n_15465 =  x_2356 & ~n_15462;
assign n_15466 = ~n_15461 &  n_15465;
assign n_15467 =  n_14817 & ~n_15466;
assign n_15468 = ~n_15464 &  n_15467;
assign n_15469 =  x_756 & ~n_14810;
assign n_15470 = ~x_1908 &  n_15440;
assign n_15471 =  x_1908 & ~n_15440;
assign n_15472 = ~n_15470 & ~n_15471;
assign n_15473 = ~n_15444 & ~n_15448;
assign n_15474 =  n_15472 & ~n_15473;
assign n_15475 = ~n_15472 &  n_15473;
assign n_15476 = ~n_15474 & ~n_15475;
assign n_15477 = ~x_692 & ~n_15476;
assign n_15478 =  x_692 & ~n_15475;
assign n_15479 = ~n_15474 &  n_15478;
assign n_15480 =  n_14812 & ~n_15479;
assign n_15481 = ~n_15477 &  n_15480;
assign n_15482 = ~n_15469 & ~n_15481;
assign n_15483 = ~n_15468 &  n_15482;
assign n_15484 =  x_756 & ~n_15483;
assign n_15485 = ~x_756 &  n_15483;
assign n_15486 = ~n_15484 & ~n_15485;
assign n_15487 = ~x_2643 &  n_15457;
assign n_15488 =  x_2643 & ~n_15457;
assign n_15489 = ~n_15487 & ~n_15488;
assign n_15490 = ~n_15461 & ~n_15465;
assign n_15491 =  n_15489 & ~n_15490;
assign n_15492 = ~n_15489 &  n_15490;
assign n_15493 = ~n_15491 & ~n_15492;
assign n_15494 = ~x_2355 & ~n_15493;
assign n_15495 =  x_2355 & ~n_15492;
assign n_15496 = ~n_15491 &  n_15495;
assign n_15497 =  n_14817 & ~n_15496;
assign n_15498 = ~n_15494 &  n_15497;
assign n_15499 =  x_755 & ~n_14810;
assign n_15500 = ~x_1907 &  n_15470;
assign n_15501 =  x_1907 & ~n_15470;
assign n_15502 = ~n_15500 & ~n_15501;
assign n_15503 = ~n_15474 & ~n_15478;
assign n_15504 =  n_15502 & ~n_15503;
assign n_15505 = ~n_15502 &  n_15503;
assign n_15506 = ~n_15504 & ~n_15505;
assign n_15507 = ~x_691 & ~n_15506;
assign n_15508 =  x_691 & ~n_15505;
assign n_15509 = ~n_15504 &  n_15508;
assign n_15510 =  n_14812 & ~n_15509;
assign n_15511 = ~n_15507 &  n_15510;
assign n_15512 = ~n_15499 & ~n_15511;
assign n_15513 = ~n_15498 &  n_15512;
assign n_15514 =  x_755 & ~n_15513;
assign n_15515 = ~x_755 &  n_15513;
assign n_15516 = ~n_15514 & ~n_15515;
assign n_15517 = ~x_2642 &  n_15487;
assign n_15518 =  x_2642 & ~n_15487;
assign n_15519 = ~n_15517 & ~n_15518;
assign n_15520 = ~n_15491 & ~n_15495;
assign n_15521 =  n_15519 & ~n_15520;
assign n_15522 = ~n_15519 &  n_15520;
assign n_15523 = ~n_15521 & ~n_15522;
assign n_15524 = ~x_2354 & ~n_15523;
assign n_15525 =  x_2354 & ~n_15522;
assign n_15526 = ~n_15521 &  n_15525;
assign n_15527 =  n_14817 & ~n_15526;
assign n_15528 = ~n_15524 &  n_15527;
assign n_15529 =  x_754 & ~n_14810;
assign n_15530 = ~x_1906 &  n_15500;
assign n_15531 =  x_1906 & ~n_15500;
assign n_15532 = ~n_15530 & ~n_15531;
assign n_15533 = ~n_15504 & ~n_15508;
assign n_15534 =  n_15532 & ~n_15533;
assign n_15535 = ~n_15532 &  n_15533;
assign n_15536 = ~n_15534 & ~n_15535;
assign n_15537 = ~x_690 & ~n_15536;
assign n_15538 =  x_690 & ~n_15535;
assign n_15539 = ~n_15534 &  n_15538;
assign n_15540 =  n_14812 & ~n_15539;
assign n_15541 = ~n_15537 &  n_15540;
assign n_15542 = ~n_15529 & ~n_15541;
assign n_15543 = ~n_15528 &  n_15542;
assign n_15544 =  x_754 & ~n_15543;
assign n_15545 = ~x_754 &  n_15543;
assign n_15546 = ~n_15544 & ~n_15545;
assign n_15547 = ~x_2641 &  n_15517;
assign n_15548 =  x_2641 & ~n_15517;
assign n_15549 = ~n_15547 & ~n_15548;
assign n_15550 = ~n_15521 & ~n_15525;
assign n_15551 =  n_15549 & ~n_15550;
assign n_15552 = ~n_15549 &  n_15550;
assign n_15553 = ~n_15551 & ~n_15552;
assign n_15554 = ~x_2353 & ~n_15553;
assign n_15555 =  x_2353 & ~n_15552;
assign n_15556 = ~n_15551 &  n_15555;
assign n_15557 =  n_14817 & ~n_15556;
assign n_15558 = ~n_15554 &  n_15557;
assign n_15559 =  x_753 & ~n_14810;
assign n_15560 = ~x_1905 &  n_15530;
assign n_15561 =  x_1905 & ~n_15530;
assign n_15562 = ~n_15560 & ~n_15561;
assign n_15563 = ~n_15534 & ~n_15538;
assign n_15564 =  n_15562 & ~n_15563;
assign n_15565 = ~n_15562 &  n_15563;
assign n_15566 = ~n_15564 & ~n_15565;
assign n_15567 = ~x_689 & ~n_15566;
assign n_15568 =  x_689 & ~n_15565;
assign n_15569 = ~n_15564 &  n_15568;
assign n_15570 =  n_14812 & ~n_15569;
assign n_15571 = ~n_15567 &  n_15570;
assign n_15572 = ~n_15559 & ~n_15571;
assign n_15573 = ~n_15558 &  n_15572;
assign n_15574 =  x_753 & ~n_15573;
assign n_15575 = ~x_753 &  n_15573;
assign n_15576 = ~n_15574 & ~n_15575;
assign n_15577 = ~x_2640 &  n_15547;
assign n_15578 =  x_2640 & ~n_15547;
assign n_15579 = ~n_15577 & ~n_15578;
assign n_15580 = ~n_15551 & ~n_15555;
assign n_15581 =  n_15579 & ~n_15580;
assign n_15582 = ~n_15579 &  n_15580;
assign n_15583 = ~n_15581 & ~n_15582;
assign n_15584 = ~x_2352 & ~n_15583;
assign n_15585 =  x_2352 & ~n_15582;
assign n_15586 = ~n_15581 &  n_15585;
assign n_15587 =  n_14817 & ~n_15586;
assign n_15588 = ~n_15584 &  n_15587;
assign n_15589 =  x_752 & ~n_14810;
assign n_15590 = ~x_1904 &  n_15560;
assign n_15591 =  x_1904 & ~n_15560;
assign n_15592 = ~n_15590 & ~n_15591;
assign n_15593 = ~n_15564 & ~n_15568;
assign n_15594 =  n_15592 & ~n_15593;
assign n_15595 = ~n_15592 &  n_15593;
assign n_15596 = ~n_15594 & ~n_15595;
assign n_15597 = ~x_688 & ~n_15596;
assign n_15598 =  x_688 & ~n_15595;
assign n_15599 = ~n_15594 &  n_15598;
assign n_15600 =  n_14812 & ~n_15599;
assign n_15601 = ~n_15597 &  n_15600;
assign n_15602 = ~n_15589 & ~n_15601;
assign n_15603 = ~n_15588 &  n_15602;
assign n_15604 =  x_752 & ~n_15603;
assign n_15605 = ~x_752 &  n_15603;
assign n_15606 = ~n_15604 & ~n_15605;
assign n_15607 = ~x_2639 &  n_15577;
assign n_15608 =  x_2639 & ~n_15577;
assign n_15609 = ~n_15607 & ~n_15608;
assign n_15610 = ~n_15581 & ~n_15585;
assign n_15611 =  n_15609 & ~n_15610;
assign n_15612 = ~n_15609 &  n_15610;
assign n_15613 = ~n_15611 & ~n_15612;
assign n_15614 = ~x_2351 & ~n_15613;
assign n_15615 =  x_2351 & ~n_15612;
assign n_15616 = ~n_15611 &  n_15615;
assign n_15617 =  n_14817 & ~n_15616;
assign n_15618 = ~n_15614 &  n_15617;
assign n_15619 =  x_751 & ~n_14810;
assign n_15620 = ~x_1903 &  n_15590;
assign n_15621 =  x_1903 & ~n_15590;
assign n_15622 = ~n_15620 & ~n_15621;
assign n_15623 = ~n_15594 & ~n_15598;
assign n_15624 =  n_15622 & ~n_15623;
assign n_15625 = ~n_15622 &  n_15623;
assign n_15626 = ~n_15624 & ~n_15625;
assign n_15627 = ~x_687 & ~n_15626;
assign n_15628 =  x_687 & ~n_15625;
assign n_15629 = ~n_15624 &  n_15628;
assign n_15630 =  n_14812 & ~n_15629;
assign n_15631 = ~n_15627 &  n_15630;
assign n_15632 = ~n_15619 & ~n_15631;
assign n_15633 = ~n_15618 &  n_15632;
assign n_15634 =  x_751 & ~n_15633;
assign n_15635 = ~x_751 &  n_15633;
assign n_15636 = ~n_15634 & ~n_15635;
assign n_15637 = ~x_2638 &  n_15607;
assign n_15638 =  x_2638 & ~n_15607;
assign n_15639 = ~n_15637 & ~n_15638;
assign n_15640 = ~n_15611 & ~n_15615;
assign n_15641 =  n_15639 & ~n_15640;
assign n_15642 = ~n_15639 &  n_15640;
assign n_15643 = ~n_15641 & ~n_15642;
assign n_15644 = ~x_2350 & ~n_15643;
assign n_15645 =  x_2350 & ~n_15642;
assign n_15646 = ~n_15641 &  n_15645;
assign n_15647 =  n_14817 & ~n_15646;
assign n_15648 = ~n_15644 &  n_15647;
assign n_15649 =  x_750 & ~n_14810;
assign n_15650 = ~x_1902 &  n_15620;
assign n_15651 =  x_1902 & ~n_15620;
assign n_15652 = ~n_15650 & ~n_15651;
assign n_15653 = ~n_15624 & ~n_15628;
assign n_15654 =  n_15652 & ~n_15653;
assign n_15655 = ~n_15652 &  n_15653;
assign n_15656 = ~n_15654 & ~n_15655;
assign n_15657 = ~x_686 & ~n_15656;
assign n_15658 =  x_686 & ~n_15655;
assign n_15659 = ~n_15654 &  n_15658;
assign n_15660 =  n_14812 & ~n_15659;
assign n_15661 = ~n_15657 &  n_15660;
assign n_15662 = ~n_15649 & ~n_15661;
assign n_15663 = ~n_15648 &  n_15662;
assign n_15664 =  x_750 & ~n_15663;
assign n_15665 = ~x_750 &  n_15663;
assign n_15666 = ~n_15664 & ~n_15665;
assign n_15667 = ~x_2637 &  n_15637;
assign n_15668 =  x_2637 & ~n_15637;
assign n_15669 = ~n_15667 & ~n_15668;
assign n_15670 = ~n_15641 & ~n_15645;
assign n_15671 =  n_15669 & ~n_15670;
assign n_15672 = ~n_15669 &  n_15670;
assign n_15673 = ~n_15671 & ~n_15672;
assign n_15674 = ~x_2349 & ~n_15673;
assign n_15675 =  x_2349 & ~n_15672;
assign n_15676 = ~n_15671 &  n_15675;
assign n_15677 =  n_14817 & ~n_15676;
assign n_15678 = ~n_15674 &  n_15677;
assign n_15679 =  x_749 & ~n_14810;
assign n_15680 = ~x_1901 &  n_15650;
assign n_15681 =  x_1901 & ~n_15650;
assign n_15682 = ~n_15680 & ~n_15681;
assign n_15683 = ~n_15654 & ~n_15658;
assign n_15684 =  n_15682 & ~n_15683;
assign n_15685 = ~n_15682 &  n_15683;
assign n_15686 = ~n_15684 & ~n_15685;
assign n_15687 = ~x_685 & ~n_15686;
assign n_15688 =  x_685 & ~n_15685;
assign n_15689 = ~n_15684 &  n_15688;
assign n_15690 =  n_14812 & ~n_15689;
assign n_15691 = ~n_15687 &  n_15690;
assign n_15692 = ~n_15679 & ~n_15691;
assign n_15693 = ~n_15678 &  n_15692;
assign n_15694 =  x_749 & ~n_15693;
assign n_15695 = ~x_749 &  n_15693;
assign n_15696 = ~n_15694 & ~n_15695;
assign n_15697 = ~x_2636 &  n_15667;
assign n_15698 =  x_2636 & ~n_15667;
assign n_15699 = ~n_15697 & ~n_15698;
assign n_15700 = ~n_15671 & ~n_15675;
assign n_15701 =  n_15699 & ~n_15700;
assign n_15702 = ~n_15699 &  n_15700;
assign n_15703 = ~n_15701 & ~n_15702;
assign n_15704 = ~x_2348 & ~n_15703;
assign n_15705 =  x_2348 & ~n_15702;
assign n_15706 = ~n_15701 &  n_15705;
assign n_15707 =  n_14817 & ~n_15706;
assign n_15708 = ~n_15704 &  n_15707;
assign n_15709 =  x_748 & ~n_14810;
assign n_15710 = ~x_1900 &  n_15680;
assign n_15711 =  x_1900 & ~n_15680;
assign n_15712 = ~n_15710 & ~n_15711;
assign n_15713 = ~n_15684 & ~n_15688;
assign n_15714 =  n_15712 & ~n_15713;
assign n_15715 = ~n_15712 &  n_15713;
assign n_15716 = ~n_15714 & ~n_15715;
assign n_15717 = ~x_684 & ~n_15716;
assign n_15718 =  x_684 & ~n_15715;
assign n_15719 = ~n_15714 &  n_15718;
assign n_15720 =  n_14812 & ~n_15719;
assign n_15721 = ~n_15717 &  n_15720;
assign n_15722 = ~n_15709 & ~n_15721;
assign n_15723 = ~n_15708 &  n_15722;
assign n_15724 =  x_748 & ~n_15723;
assign n_15725 = ~x_748 &  n_15723;
assign n_15726 = ~n_15724 & ~n_15725;
assign n_15727 = ~n_15714 & ~n_15718;
assign n_15728 =  x_683 & ~x_1899;
assign n_15729 = ~x_683 &  x_1899;
assign n_15730 = ~n_15728 & ~n_15729;
assign n_15731 =  n_15710 &  n_15730;
assign n_15732 = ~n_15710 & ~n_15730;
assign n_15733 = ~n_15731 & ~n_15732;
assign n_15734 =  n_15727 & ~n_15733;
assign n_15735 = ~n_15727 &  n_15733;
assign n_15736 =  n_14812 & ~n_15735;
assign n_15737 = ~n_15734 &  n_15736;
assign n_15738 =  x_747 & ~n_14810;
assign n_15739 = ~n_15701 & ~n_15705;
assign n_15740 =  x_2347 & ~x_2635;
assign n_15741 = ~x_2347 &  x_2635;
assign n_15742 = ~n_15740 & ~n_15741;
assign n_15743 =  n_15697 &  n_15742;
assign n_15744 = ~n_15697 & ~n_15742;
assign n_15745 = ~n_15743 & ~n_15744;
assign n_15746 =  n_15739 & ~n_15745;
assign n_15747 = ~n_15739 &  n_15745;
assign n_15748 =  n_14817 & ~n_15747;
assign n_15749 = ~n_15746 &  n_15748;
assign n_15750 = ~n_15738 & ~n_15749;
assign n_15751 = ~n_15737 &  n_15750;
assign n_15752 =  x_747 & ~n_15751;
assign n_15753 = ~x_747 &  n_15751;
assign n_15754 = ~n_15752 & ~n_15753;
assign n_15755 =  n_12614 &  n_6331;
assign n_15756 =  x_746 & ~n_15755;
assign n_15757 =  i_32 &  n_15755;
assign n_15758 = ~n_15756 & ~n_15757;
assign n_15759 =  x_746 & ~n_15758;
assign n_15760 = ~x_746 &  n_15758;
assign n_15761 = ~n_15759 & ~n_15760;
assign n_15762 =  x_745 & ~n_15755;
assign n_15763 =  i_31 &  n_15755;
assign n_15764 = ~n_15762 & ~n_15763;
assign n_15765 =  x_745 & ~n_15764;
assign n_15766 = ~x_745 &  n_15764;
assign n_15767 = ~n_15765 & ~n_15766;
assign n_15768 =  x_744 & ~n_15755;
assign n_15769 =  i_30 &  n_15755;
assign n_15770 = ~n_15768 & ~n_15769;
assign n_15771 =  x_744 & ~n_15770;
assign n_15772 = ~x_744 &  n_15770;
assign n_15773 = ~n_15771 & ~n_15772;
assign n_15774 =  x_743 & ~n_15755;
assign n_15775 =  i_29 &  n_15755;
assign n_15776 = ~n_15774 & ~n_15775;
assign n_15777 =  x_743 & ~n_15776;
assign n_15778 = ~x_743 &  n_15776;
assign n_15779 = ~n_15777 & ~n_15778;
assign n_15780 =  x_742 & ~n_15755;
assign n_15781 =  i_28 &  n_15755;
assign n_15782 = ~n_15780 & ~n_15781;
assign n_15783 =  x_742 & ~n_15782;
assign n_15784 = ~x_742 &  n_15782;
assign n_15785 = ~n_15783 & ~n_15784;
assign n_15786 =  x_741 & ~n_15755;
assign n_15787 =  i_27 &  n_15755;
assign n_15788 = ~n_15786 & ~n_15787;
assign n_15789 =  x_741 & ~n_15788;
assign n_15790 = ~x_741 &  n_15788;
assign n_15791 = ~n_15789 & ~n_15790;
assign n_15792 =  x_740 & ~n_15755;
assign n_15793 =  i_26 &  n_15755;
assign n_15794 = ~n_15792 & ~n_15793;
assign n_15795 =  x_740 & ~n_15794;
assign n_15796 = ~x_740 &  n_15794;
assign n_15797 = ~n_15795 & ~n_15796;
assign n_15798 =  x_739 & ~n_15755;
assign n_15799 =  i_25 &  n_15755;
assign n_15800 = ~n_15798 & ~n_15799;
assign n_15801 =  x_739 & ~n_15800;
assign n_15802 = ~x_739 &  n_15800;
assign n_15803 = ~n_15801 & ~n_15802;
assign n_15804 =  x_738 & ~n_15755;
assign n_15805 =  i_24 &  n_15755;
assign n_15806 = ~n_15804 & ~n_15805;
assign n_15807 =  x_738 & ~n_15806;
assign n_15808 = ~x_738 &  n_15806;
assign n_15809 = ~n_15807 & ~n_15808;
assign n_15810 =  x_737 & ~n_15755;
assign n_15811 =  i_23 &  n_15755;
assign n_15812 = ~n_15810 & ~n_15811;
assign n_15813 =  x_737 & ~n_15812;
assign n_15814 = ~x_737 &  n_15812;
assign n_15815 = ~n_15813 & ~n_15814;
assign n_15816 =  x_736 & ~n_15755;
assign n_15817 =  i_22 &  n_15755;
assign n_15818 = ~n_15816 & ~n_15817;
assign n_15819 =  x_736 & ~n_15818;
assign n_15820 = ~x_736 &  n_15818;
assign n_15821 = ~n_15819 & ~n_15820;
assign n_15822 =  x_735 & ~n_15755;
assign n_15823 =  i_21 &  n_15755;
assign n_15824 = ~n_15822 & ~n_15823;
assign n_15825 =  x_735 & ~n_15824;
assign n_15826 = ~x_735 &  n_15824;
assign n_15827 = ~n_15825 & ~n_15826;
assign n_15828 =  x_734 & ~n_15755;
assign n_15829 =  i_20 &  n_15755;
assign n_15830 = ~n_15828 & ~n_15829;
assign n_15831 =  x_734 & ~n_15830;
assign n_15832 = ~x_734 &  n_15830;
assign n_15833 = ~n_15831 & ~n_15832;
assign n_15834 =  x_733 & ~n_15755;
assign n_15835 =  i_19 &  n_15755;
assign n_15836 = ~n_15834 & ~n_15835;
assign n_15837 =  x_733 & ~n_15836;
assign n_15838 = ~x_733 &  n_15836;
assign n_15839 = ~n_15837 & ~n_15838;
assign n_15840 =  x_732 & ~n_15755;
assign n_15841 =  i_18 &  n_15755;
assign n_15842 = ~n_15840 & ~n_15841;
assign n_15843 =  x_732 & ~n_15842;
assign n_15844 = ~x_732 &  n_15842;
assign n_15845 = ~n_15843 & ~n_15844;
assign n_15846 =  x_731 & ~n_15755;
assign n_15847 =  i_17 &  n_15755;
assign n_15848 = ~n_15846 & ~n_15847;
assign n_15849 =  x_731 & ~n_15848;
assign n_15850 = ~x_731 &  n_15848;
assign n_15851 = ~n_15849 & ~n_15850;
assign n_15852 =  x_730 & ~n_15755;
assign n_15853 =  i_16 &  n_15755;
assign n_15854 = ~n_15852 & ~n_15853;
assign n_15855 =  x_730 & ~n_15854;
assign n_15856 = ~x_730 &  n_15854;
assign n_15857 = ~n_15855 & ~n_15856;
assign n_15858 =  x_729 & ~n_15755;
assign n_15859 =  i_15 &  n_15755;
assign n_15860 = ~n_15858 & ~n_15859;
assign n_15861 =  x_729 & ~n_15860;
assign n_15862 = ~x_729 &  n_15860;
assign n_15863 = ~n_15861 & ~n_15862;
assign n_15864 =  x_728 & ~n_15755;
assign n_15865 =  i_14 &  n_15755;
assign n_15866 = ~n_15864 & ~n_15865;
assign n_15867 =  x_728 & ~n_15866;
assign n_15868 = ~x_728 &  n_15866;
assign n_15869 = ~n_15867 & ~n_15868;
assign n_15870 =  x_727 & ~n_15755;
assign n_15871 =  i_13 &  n_15755;
assign n_15872 = ~n_15870 & ~n_15871;
assign n_15873 =  x_727 & ~n_15872;
assign n_15874 = ~x_727 &  n_15872;
assign n_15875 = ~n_15873 & ~n_15874;
assign n_15876 =  x_726 & ~n_15755;
assign n_15877 =  i_12 &  n_15755;
assign n_15878 = ~n_15876 & ~n_15877;
assign n_15879 =  x_726 & ~n_15878;
assign n_15880 = ~x_726 &  n_15878;
assign n_15881 = ~n_15879 & ~n_15880;
assign n_15882 =  x_725 & ~n_15755;
assign n_15883 =  i_11 &  n_15755;
assign n_15884 = ~n_15882 & ~n_15883;
assign n_15885 =  x_725 & ~n_15884;
assign n_15886 = ~x_725 &  n_15884;
assign n_15887 = ~n_15885 & ~n_15886;
assign n_15888 =  x_724 & ~n_15755;
assign n_15889 =  i_10 &  n_15755;
assign n_15890 = ~n_15888 & ~n_15889;
assign n_15891 =  x_724 & ~n_15890;
assign n_15892 = ~x_724 &  n_15890;
assign n_15893 = ~n_15891 & ~n_15892;
assign n_15894 =  x_723 & ~n_15755;
assign n_15895 =  i_9 &  n_15755;
assign n_15896 = ~n_15894 & ~n_15895;
assign n_15897 =  x_723 & ~n_15896;
assign n_15898 = ~x_723 &  n_15896;
assign n_15899 = ~n_15897 & ~n_15898;
assign n_15900 =  x_722 & ~n_15755;
assign n_15901 =  i_8 &  n_15755;
assign n_15902 = ~n_15900 & ~n_15901;
assign n_15903 =  x_722 & ~n_15902;
assign n_15904 = ~x_722 &  n_15902;
assign n_15905 = ~n_15903 & ~n_15904;
assign n_15906 =  x_721 & ~n_15755;
assign n_15907 =  i_7 &  n_15755;
assign n_15908 = ~n_15906 & ~n_15907;
assign n_15909 =  x_721 & ~n_15908;
assign n_15910 = ~x_721 &  n_15908;
assign n_15911 = ~n_15909 & ~n_15910;
assign n_15912 =  x_720 & ~n_15755;
assign n_15913 =  i_6 &  n_15755;
assign n_15914 = ~n_15912 & ~n_15913;
assign n_15915 =  x_720 & ~n_15914;
assign n_15916 = ~x_720 &  n_15914;
assign n_15917 = ~n_15915 & ~n_15916;
assign n_15918 =  x_719 & ~n_15755;
assign n_15919 =  i_5 &  n_15755;
assign n_15920 = ~n_15918 & ~n_15919;
assign n_15921 =  x_719 & ~n_15920;
assign n_15922 = ~x_719 &  n_15920;
assign n_15923 = ~n_15921 & ~n_15922;
assign n_15924 =  x_718 & ~n_15755;
assign n_15925 =  i_4 &  n_15755;
assign n_15926 = ~n_15924 & ~n_15925;
assign n_15927 =  x_718 & ~n_15926;
assign n_15928 = ~x_718 &  n_15926;
assign n_15929 = ~n_15927 & ~n_15928;
assign n_15930 =  x_717 & ~n_15755;
assign n_15931 =  i_3 &  n_15755;
assign n_15932 = ~n_15930 & ~n_15931;
assign n_15933 =  x_717 & ~n_15932;
assign n_15934 = ~x_717 &  n_15932;
assign n_15935 = ~n_15933 & ~n_15934;
assign n_15936 =  x_716 & ~n_15755;
assign n_15937 =  i_2 &  n_15755;
assign n_15938 = ~n_15936 & ~n_15937;
assign n_15939 =  x_716 & ~n_15938;
assign n_15940 = ~x_716 &  n_15938;
assign n_15941 = ~n_15939 & ~n_15940;
assign n_15942 =  x_715 & ~n_15755;
assign n_15943 =  i_1 &  n_15755;
assign n_15944 = ~n_15942 & ~n_15943;
assign n_15945 =  x_715 & ~n_15944;
assign n_15946 = ~x_715 &  n_15944;
assign n_15947 = ~n_15945 & ~n_15946;
assign n_15948 =  n_4993 &  n_8;
assign n_15949 =  x_714 & ~n_15948;
assign n_15950 =  i_32 &  n_15948;
assign n_15951 = ~n_15949 & ~n_15950;
assign n_15952 =  x_714 & ~n_15951;
assign n_15953 = ~x_714 &  n_15951;
assign n_15954 = ~n_15952 & ~n_15953;
assign n_15955 =  x_713 & ~n_15948;
assign n_15956 =  i_31 &  n_15948;
assign n_15957 = ~n_15955 & ~n_15956;
assign n_15958 =  x_713 & ~n_15957;
assign n_15959 = ~x_713 &  n_15957;
assign n_15960 = ~n_15958 & ~n_15959;
assign n_15961 =  x_712 & ~n_15948;
assign n_15962 =  i_30 &  n_15948;
assign n_15963 = ~n_15961 & ~n_15962;
assign n_15964 =  x_712 & ~n_15963;
assign n_15965 = ~x_712 &  n_15963;
assign n_15966 = ~n_15964 & ~n_15965;
assign n_15967 =  x_711 & ~n_15948;
assign n_15968 =  i_29 &  n_15948;
assign n_15969 = ~n_15967 & ~n_15968;
assign n_15970 =  x_711 & ~n_15969;
assign n_15971 = ~x_711 &  n_15969;
assign n_15972 = ~n_15970 & ~n_15971;
assign n_15973 =  x_710 & ~n_15948;
assign n_15974 =  i_28 &  n_15948;
assign n_15975 = ~n_15973 & ~n_15974;
assign n_15976 =  x_710 & ~n_15975;
assign n_15977 = ~x_710 &  n_15975;
assign n_15978 = ~n_15976 & ~n_15977;
assign n_15979 =  x_709 & ~n_15948;
assign n_15980 =  i_27 &  n_15948;
assign n_15981 = ~n_15979 & ~n_15980;
assign n_15982 =  x_709 & ~n_15981;
assign n_15983 = ~x_709 &  n_15981;
assign n_15984 = ~n_15982 & ~n_15983;
assign n_15985 =  x_708 & ~n_15948;
assign n_15986 =  i_26 &  n_15948;
assign n_15987 = ~n_15985 & ~n_15986;
assign n_15988 =  x_708 & ~n_15987;
assign n_15989 = ~x_708 &  n_15987;
assign n_15990 = ~n_15988 & ~n_15989;
assign n_15991 =  x_707 & ~n_15948;
assign n_15992 =  i_25 &  n_15948;
assign n_15993 = ~n_15991 & ~n_15992;
assign n_15994 =  x_707 & ~n_15993;
assign n_15995 = ~x_707 &  n_15993;
assign n_15996 = ~n_15994 & ~n_15995;
assign n_15997 =  x_706 & ~n_15948;
assign n_15998 =  i_24 &  n_15948;
assign n_15999 = ~n_15997 & ~n_15998;
assign n_16000 =  x_706 & ~n_15999;
assign n_16001 = ~x_706 &  n_15999;
assign n_16002 = ~n_16000 & ~n_16001;
assign n_16003 =  x_705 & ~n_15948;
assign n_16004 =  i_23 &  n_15948;
assign n_16005 = ~n_16003 & ~n_16004;
assign n_16006 =  x_705 & ~n_16005;
assign n_16007 = ~x_705 &  n_16005;
assign n_16008 = ~n_16006 & ~n_16007;
assign n_16009 =  x_704 & ~n_15948;
assign n_16010 =  i_22 &  n_15948;
assign n_16011 = ~n_16009 & ~n_16010;
assign n_16012 =  x_704 & ~n_16011;
assign n_16013 = ~x_704 &  n_16011;
assign n_16014 = ~n_16012 & ~n_16013;
assign n_16015 =  x_703 & ~n_15948;
assign n_16016 =  i_21 &  n_15948;
assign n_16017 = ~n_16015 & ~n_16016;
assign n_16018 =  x_703 & ~n_16017;
assign n_16019 = ~x_703 &  n_16017;
assign n_16020 = ~n_16018 & ~n_16019;
assign n_16021 =  x_702 & ~n_15948;
assign n_16022 =  i_20 &  n_15948;
assign n_16023 = ~n_16021 & ~n_16022;
assign n_16024 =  x_702 & ~n_16023;
assign n_16025 = ~x_702 &  n_16023;
assign n_16026 = ~n_16024 & ~n_16025;
assign n_16027 =  x_701 & ~n_15948;
assign n_16028 =  i_19 &  n_15948;
assign n_16029 = ~n_16027 & ~n_16028;
assign n_16030 =  x_701 & ~n_16029;
assign n_16031 = ~x_701 &  n_16029;
assign n_16032 = ~n_16030 & ~n_16031;
assign n_16033 =  x_700 & ~n_15948;
assign n_16034 =  i_18 &  n_15948;
assign n_16035 = ~n_16033 & ~n_16034;
assign n_16036 =  x_700 & ~n_16035;
assign n_16037 = ~x_700 &  n_16035;
assign n_16038 = ~n_16036 & ~n_16037;
assign n_16039 =  x_699 & ~n_15948;
assign n_16040 =  i_17 &  n_15948;
assign n_16041 = ~n_16039 & ~n_16040;
assign n_16042 =  x_699 & ~n_16041;
assign n_16043 = ~x_699 &  n_16041;
assign n_16044 = ~n_16042 & ~n_16043;
assign n_16045 =  x_698 & ~n_15948;
assign n_16046 =  i_16 &  n_15948;
assign n_16047 = ~n_16045 & ~n_16046;
assign n_16048 =  x_698 & ~n_16047;
assign n_16049 = ~x_698 &  n_16047;
assign n_16050 = ~n_16048 & ~n_16049;
assign n_16051 =  x_697 & ~n_15948;
assign n_16052 =  i_15 &  n_15948;
assign n_16053 = ~n_16051 & ~n_16052;
assign n_16054 =  x_697 & ~n_16053;
assign n_16055 = ~x_697 &  n_16053;
assign n_16056 = ~n_16054 & ~n_16055;
assign n_16057 =  x_696 & ~n_15948;
assign n_16058 =  i_14 &  n_15948;
assign n_16059 = ~n_16057 & ~n_16058;
assign n_16060 =  x_696 & ~n_16059;
assign n_16061 = ~x_696 &  n_16059;
assign n_16062 = ~n_16060 & ~n_16061;
assign n_16063 =  x_695 & ~n_15948;
assign n_16064 =  i_13 &  n_15948;
assign n_16065 = ~n_16063 & ~n_16064;
assign n_16066 =  x_695 & ~n_16065;
assign n_16067 = ~x_695 &  n_16065;
assign n_16068 = ~n_16066 & ~n_16067;
assign n_16069 =  x_694 & ~n_15948;
assign n_16070 =  i_12 &  n_15948;
assign n_16071 = ~n_16069 & ~n_16070;
assign n_16072 =  x_694 & ~n_16071;
assign n_16073 = ~x_694 &  n_16071;
assign n_16074 = ~n_16072 & ~n_16073;
assign n_16075 =  x_693 & ~n_15948;
assign n_16076 =  i_11 &  n_15948;
assign n_16077 = ~n_16075 & ~n_16076;
assign n_16078 =  x_693 & ~n_16077;
assign n_16079 = ~x_693 &  n_16077;
assign n_16080 = ~n_16078 & ~n_16079;
assign n_16081 =  x_692 & ~n_15948;
assign n_16082 =  i_10 &  n_15948;
assign n_16083 = ~n_16081 & ~n_16082;
assign n_16084 =  x_692 & ~n_16083;
assign n_16085 = ~x_692 &  n_16083;
assign n_16086 = ~n_16084 & ~n_16085;
assign n_16087 =  x_691 & ~n_15948;
assign n_16088 =  i_9 &  n_15948;
assign n_16089 = ~n_16087 & ~n_16088;
assign n_16090 =  x_691 & ~n_16089;
assign n_16091 = ~x_691 &  n_16089;
assign n_16092 = ~n_16090 & ~n_16091;
assign n_16093 =  x_690 & ~n_15948;
assign n_16094 =  i_8 &  n_15948;
assign n_16095 = ~n_16093 & ~n_16094;
assign n_16096 =  x_690 & ~n_16095;
assign n_16097 = ~x_690 &  n_16095;
assign n_16098 = ~n_16096 & ~n_16097;
assign n_16099 =  x_689 & ~n_15948;
assign n_16100 =  i_7 &  n_15948;
assign n_16101 = ~n_16099 & ~n_16100;
assign n_16102 =  x_689 & ~n_16101;
assign n_16103 = ~x_689 &  n_16101;
assign n_16104 = ~n_16102 & ~n_16103;
assign n_16105 =  x_688 & ~n_15948;
assign n_16106 =  i_6 &  n_15948;
assign n_16107 = ~n_16105 & ~n_16106;
assign n_16108 =  x_688 & ~n_16107;
assign n_16109 = ~x_688 &  n_16107;
assign n_16110 = ~n_16108 & ~n_16109;
assign n_16111 =  x_687 & ~n_15948;
assign n_16112 =  i_5 &  n_15948;
assign n_16113 = ~n_16111 & ~n_16112;
assign n_16114 =  x_687 & ~n_16113;
assign n_16115 = ~x_687 &  n_16113;
assign n_16116 = ~n_16114 & ~n_16115;
assign n_16117 =  x_686 & ~n_15948;
assign n_16118 =  i_4 &  n_15948;
assign n_16119 = ~n_16117 & ~n_16118;
assign n_16120 =  x_686 & ~n_16119;
assign n_16121 = ~x_686 &  n_16119;
assign n_16122 = ~n_16120 & ~n_16121;
assign n_16123 =  x_685 & ~n_15948;
assign n_16124 =  i_3 &  n_15948;
assign n_16125 = ~n_16123 & ~n_16124;
assign n_16126 =  x_685 & ~n_16125;
assign n_16127 = ~x_685 &  n_16125;
assign n_16128 = ~n_16126 & ~n_16127;
assign n_16129 =  x_684 & ~n_15948;
assign n_16130 =  i_2 &  n_15948;
assign n_16131 = ~n_16129 & ~n_16130;
assign n_16132 =  x_684 & ~n_16131;
assign n_16133 = ~x_684 &  n_16131;
assign n_16134 = ~n_16132 & ~n_16133;
assign n_16135 =  x_683 & ~n_15948;
assign n_16136 =  i_1 &  n_15948;
assign n_16137 = ~n_16135 & ~n_16136;
assign n_16138 =  x_683 & ~n_16137;
assign n_16139 = ~x_683 &  n_16137;
assign n_16140 = ~n_16138 & ~n_16139;
assign n_16141 =  n_4993 &  n_2101;
assign n_16142 =  x_682 & ~n_16141;
assign n_16143 =  i_32 &  n_16141;
assign n_16144 = ~n_16142 & ~n_16143;
assign n_16145 =  x_682 & ~n_16144;
assign n_16146 = ~x_682 &  n_16144;
assign n_16147 = ~n_16145 & ~n_16146;
assign n_16148 =  x_681 & ~n_16141;
assign n_16149 =  i_31 &  n_16141;
assign n_16150 = ~n_16148 & ~n_16149;
assign n_16151 =  x_681 & ~n_16150;
assign n_16152 = ~x_681 &  n_16150;
assign n_16153 = ~n_16151 & ~n_16152;
assign n_16154 =  x_680 & ~n_16141;
assign n_16155 =  i_30 &  n_16141;
assign n_16156 = ~n_16154 & ~n_16155;
assign n_16157 =  x_680 & ~n_16156;
assign n_16158 = ~x_680 &  n_16156;
assign n_16159 = ~n_16157 & ~n_16158;
assign n_16160 =  x_679 & ~n_16141;
assign n_16161 =  i_29 &  n_16141;
assign n_16162 = ~n_16160 & ~n_16161;
assign n_16163 =  x_679 & ~n_16162;
assign n_16164 = ~x_679 &  n_16162;
assign n_16165 = ~n_16163 & ~n_16164;
assign n_16166 =  x_678 & ~n_16141;
assign n_16167 =  i_28 &  n_16141;
assign n_16168 = ~n_16166 & ~n_16167;
assign n_16169 =  x_678 & ~n_16168;
assign n_16170 = ~x_678 &  n_16168;
assign n_16171 = ~n_16169 & ~n_16170;
assign n_16172 =  x_677 & ~n_16141;
assign n_16173 =  i_27 &  n_16141;
assign n_16174 = ~n_16172 & ~n_16173;
assign n_16175 =  x_677 & ~n_16174;
assign n_16176 = ~x_677 &  n_16174;
assign n_16177 = ~n_16175 & ~n_16176;
assign n_16178 =  x_676 & ~n_16141;
assign n_16179 =  i_26 &  n_16141;
assign n_16180 = ~n_16178 & ~n_16179;
assign n_16181 =  x_676 & ~n_16180;
assign n_16182 = ~x_676 &  n_16180;
assign n_16183 = ~n_16181 & ~n_16182;
assign n_16184 =  x_675 & ~n_16141;
assign n_16185 =  i_25 &  n_16141;
assign n_16186 = ~n_16184 & ~n_16185;
assign n_16187 =  x_675 & ~n_16186;
assign n_16188 = ~x_675 &  n_16186;
assign n_16189 = ~n_16187 & ~n_16188;
assign n_16190 =  x_674 & ~n_16141;
assign n_16191 =  i_24 &  n_16141;
assign n_16192 = ~n_16190 & ~n_16191;
assign n_16193 =  x_674 & ~n_16192;
assign n_16194 = ~x_674 &  n_16192;
assign n_16195 = ~n_16193 & ~n_16194;
assign n_16196 =  x_673 & ~n_16141;
assign n_16197 =  i_23 &  n_16141;
assign n_16198 = ~n_16196 & ~n_16197;
assign n_16199 =  x_673 & ~n_16198;
assign n_16200 = ~x_673 &  n_16198;
assign n_16201 = ~n_16199 & ~n_16200;
assign n_16202 =  x_672 & ~n_16141;
assign n_16203 =  i_22 &  n_16141;
assign n_16204 = ~n_16202 & ~n_16203;
assign n_16205 =  x_672 & ~n_16204;
assign n_16206 = ~x_672 &  n_16204;
assign n_16207 = ~n_16205 & ~n_16206;
assign n_16208 =  x_671 & ~n_16141;
assign n_16209 =  i_21 &  n_16141;
assign n_16210 = ~n_16208 & ~n_16209;
assign n_16211 =  x_671 & ~n_16210;
assign n_16212 = ~x_671 &  n_16210;
assign n_16213 = ~n_16211 & ~n_16212;
assign n_16214 =  x_670 & ~n_16141;
assign n_16215 =  i_20 &  n_16141;
assign n_16216 = ~n_16214 & ~n_16215;
assign n_16217 =  x_670 & ~n_16216;
assign n_16218 = ~x_670 &  n_16216;
assign n_16219 = ~n_16217 & ~n_16218;
assign n_16220 =  x_669 & ~n_16141;
assign n_16221 =  i_19 &  n_16141;
assign n_16222 = ~n_16220 & ~n_16221;
assign n_16223 =  x_669 & ~n_16222;
assign n_16224 = ~x_669 &  n_16222;
assign n_16225 = ~n_16223 & ~n_16224;
assign n_16226 =  x_668 & ~n_16141;
assign n_16227 =  i_18 &  n_16141;
assign n_16228 = ~n_16226 & ~n_16227;
assign n_16229 =  x_668 & ~n_16228;
assign n_16230 = ~x_668 &  n_16228;
assign n_16231 = ~n_16229 & ~n_16230;
assign n_16232 =  x_667 & ~n_16141;
assign n_16233 =  i_17 &  n_16141;
assign n_16234 = ~n_16232 & ~n_16233;
assign n_16235 =  x_667 & ~n_16234;
assign n_16236 = ~x_667 &  n_16234;
assign n_16237 = ~n_16235 & ~n_16236;
assign n_16238 =  x_666 & ~n_16141;
assign n_16239 =  i_16 &  n_16141;
assign n_16240 = ~n_16238 & ~n_16239;
assign n_16241 =  x_666 & ~n_16240;
assign n_16242 = ~x_666 &  n_16240;
assign n_16243 = ~n_16241 & ~n_16242;
assign n_16244 =  x_665 & ~n_16141;
assign n_16245 =  i_15 &  n_16141;
assign n_16246 = ~n_16244 & ~n_16245;
assign n_16247 =  x_665 & ~n_16246;
assign n_16248 = ~x_665 &  n_16246;
assign n_16249 = ~n_16247 & ~n_16248;
assign n_16250 =  x_664 & ~n_16141;
assign n_16251 =  i_14 &  n_16141;
assign n_16252 = ~n_16250 & ~n_16251;
assign n_16253 =  x_664 & ~n_16252;
assign n_16254 = ~x_664 &  n_16252;
assign n_16255 = ~n_16253 & ~n_16254;
assign n_16256 =  x_663 & ~n_16141;
assign n_16257 =  i_13 &  n_16141;
assign n_16258 = ~n_16256 & ~n_16257;
assign n_16259 =  x_663 & ~n_16258;
assign n_16260 = ~x_663 &  n_16258;
assign n_16261 = ~n_16259 & ~n_16260;
assign n_16262 =  x_662 & ~n_16141;
assign n_16263 =  i_12 &  n_16141;
assign n_16264 = ~n_16262 & ~n_16263;
assign n_16265 =  x_662 & ~n_16264;
assign n_16266 = ~x_662 &  n_16264;
assign n_16267 = ~n_16265 & ~n_16266;
assign n_16268 =  x_661 & ~n_16141;
assign n_16269 =  i_11 &  n_16141;
assign n_16270 = ~n_16268 & ~n_16269;
assign n_16271 =  x_661 & ~n_16270;
assign n_16272 = ~x_661 &  n_16270;
assign n_16273 = ~n_16271 & ~n_16272;
assign n_16274 =  x_660 & ~n_16141;
assign n_16275 =  i_10 &  n_16141;
assign n_16276 = ~n_16274 & ~n_16275;
assign n_16277 =  x_660 & ~n_16276;
assign n_16278 = ~x_660 &  n_16276;
assign n_16279 = ~n_16277 & ~n_16278;
assign n_16280 =  x_659 & ~n_16141;
assign n_16281 =  i_9 &  n_16141;
assign n_16282 = ~n_16280 & ~n_16281;
assign n_16283 =  x_659 & ~n_16282;
assign n_16284 = ~x_659 &  n_16282;
assign n_16285 = ~n_16283 & ~n_16284;
assign n_16286 =  x_658 & ~n_16141;
assign n_16287 =  i_8 &  n_16141;
assign n_16288 = ~n_16286 & ~n_16287;
assign n_16289 =  x_658 & ~n_16288;
assign n_16290 = ~x_658 &  n_16288;
assign n_16291 = ~n_16289 & ~n_16290;
assign n_16292 =  x_657 & ~n_16141;
assign n_16293 =  i_7 &  n_16141;
assign n_16294 = ~n_16292 & ~n_16293;
assign n_16295 =  x_657 & ~n_16294;
assign n_16296 = ~x_657 &  n_16294;
assign n_16297 = ~n_16295 & ~n_16296;
assign n_16298 =  x_656 & ~n_16141;
assign n_16299 =  i_6 &  n_16141;
assign n_16300 = ~n_16298 & ~n_16299;
assign n_16301 =  x_656 & ~n_16300;
assign n_16302 = ~x_656 &  n_16300;
assign n_16303 = ~n_16301 & ~n_16302;
assign n_16304 =  x_655 & ~n_16141;
assign n_16305 =  i_5 &  n_16141;
assign n_16306 = ~n_16304 & ~n_16305;
assign n_16307 =  x_655 & ~n_16306;
assign n_16308 = ~x_655 &  n_16306;
assign n_16309 = ~n_16307 & ~n_16308;
assign n_16310 =  x_654 & ~n_16141;
assign n_16311 =  i_4 &  n_16141;
assign n_16312 = ~n_16310 & ~n_16311;
assign n_16313 =  x_654 & ~n_16312;
assign n_16314 = ~x_654 &  n_16312;
assign n_16315 = ~n_16313 & ~n_16314;
assign n_16316 =  x_653 & ~n_16141;
assign n_16317 =  i_3 &  n_16141;
assign n_16318 = ~n_16316 & ~n_16317;
assign n_16319 =  x_653 & ~n_16318;
assign n_16320 = ~x_653 &  n_16318;
assign n_16321 = ~n_16319 & ~n_16320;
assign n_16322 =  x_652 & ~n_16141;
assign n_16323 =  i_2 &  n_16141;
assign n_16324 = ~n_16322 & ~n_16323;
assign n_16325 =  x_652 & ~n_16324;
assign n_16326 = ~x_652 &  n_16324;
assign n_16327 = ~n_16325 & ~n_16326;
assign n_16328 =  x_651 & ~n_16141;
assign n_16329 =  i_1 &  n_16141;
assign n_16330 = ~n_16328 & ~n_16329;
assign n_16331 =  x_651 & ~n_16330;
assign n_16332 = ~x_651 &  n_16330;
assign n_16333 = ~n_16331 & ~n_16332;
assign n_16334 =  n_586 &  n_1904;
assign n_16335 = ~x_39 &  n_16334;
assign n_16336 =  x_650 & ~n_16335;
assign n_16337 =  i_32 &  n_16335;
assign n_16338 = ~n_16336 & ~n_16337;
assign n_16339 =  x_650 & ~n_16338;
assign n_16340 = ~x_650 &  n_16338;
assign n_16341 = ~n_16339 & ~n_16340;
assign n_16342 =  x_649 & ~n_16335;
assign n_16343 =  i_31 &  n_16335;
assign n_16344 = ~n_16342 & ~n_16343;
assign n_16345 =  x_649 & ~n_16344;
assign n_16346 = ~x_649 &  n_16344;
assign n_16347 = ~n_16345 & ~n_16346;
assign n_16348 =  x_648 & ~n_16335;
assign n_16349 =  i_30 &  n_16335;
assign n_16350 = ~n_16348 & ~n_16349;
assign n_16351 =  x_648 & ~n_16350;
assign n_16352 = ~x_648 &  n_16350;
assign n_16353 = ~n_16351 & ~n_16352;
assign n_16354 =  x_647 & ~n_16335;
assign n_16355 =  i_29 &  n_16335;
assign n_16356 = ~n_16354 & ~n_16355;
assign n_16357 =  x_647 & ~n_16356;
assign n_16358 = ~x_647 &  n_16356;
assign n_16359 = ~n_16357 & ~n_16358;
assign n_16360 =  x_646 & ~n_16335;
assign n_16361 =  i_28 &  n_16335;
assign n_16362 = ~n_16360 & ~n_16361;
assign n_16363 =  x_646 & ~n_16362;
assign n_16364 = ~x_646 &  n_16362;
assign n_16365 = ~n_16363 & ~n_16364;
assign n_16366 =  x_645 & ~n_16335;
assign n_16367 =  i_27 &  n_16335;
assign n_16368 = ~n_16366 & ~n_16367;
assign n_16369 =  x_645 & ~n_16368;
assign n_16370 = ~x_645 &  n_16368;
assign n_16371 = ~n_16369 & ~n_16370;
assign n_16372 =  x_644 & ~n_16335;
assign n_16373 =  i_26 &  n_16335;
assign n_16374 = ~n_16372 & ~n_16373;
assign n_16375 =  x_644 & ~n_16374;
assign n_16376 = ~x_644 &  n_16374;
assign n_16377 = ~n_16375 & ~n_16376;
assign n_16378 =  x_643 & ~n_16335;
assign n_16379 =  i_25 &  n_16335;
assign n_16380 = ~n_16378 & ~n_16379;
assign n_16381 =  x_643 & ~n_16380;
assign n_16382 = ~x_643 &  n_16380;
assign n_16383 = ~n_16381 & ~n_16382;
assign n_16384 =  x_642 & ~n_16335;
assign n_16385 =  i_24 &  n_16335;
assign n_16386 = ~n_16384 & ~n_16385;
assign n_16387 =  x_642 & ~n_16386;
assign n_16388 = ~x_642 &  n_16386;
assign n_16389 = ~n_16387 & ~n_16388;
assign n_16390 =  x_641 & ~n_16335;
assign n_16391 =  i_23 &  n_16335;
assign n_16392 = ~n_16390 & ~n_16391;
assign n_16393 =  x_641 & ~n_16392;
assign n_16394 = ~x_641 &  n_16392;
assign n_16395 = ~n_16393 & ~n_16394;
assign n_16396 =  x_640 & ~n_16335;
assign n_16397 =  i_22 &  n_16335;
assign n_16398 = ~n_16396 & ~n_16397;
assign n_16399 =  x_640 & ~n_16398;
assign n_16400 = ~x_640 &  n_16398;
assign n_16401 = ~n_16399 & ~n_16400;
assign n_16402 =  x_639 & ~n_16335;
assign n_16403 =  i_21 &  n_16335;
assign n_16404 = ~n_16402 & ~n_16403;
assign n_16405 =  x_639 & ~n_16404;
assign n_16406 = ~x_639 &  n_16404;
assign n_16407 = ~n_16405 & ~n_16406;
assign n_16408 =  x_638 & ~n_16335;
assign n_16409 =  i_20 &  n_16335;
assign n_16410 = ~n_16408 & ~n_16409;
assign n_16411 =  x_638 & ~n_16410;
assign n_16412 = ~x_638 &  n_16410;
assign n_16413 = ~n_16411 & ~n_16412;
assign n_16414 =  x_637 & ~n_16335;
assign n_16415 =  i_19 &  n_16335;
assign n_16416 = ~n_16414 & ~n_16415;
assign n_16417 =  x_637 & ~n_16416;
assign n_16418 = ~x_637 &  n_16416;
assign n_16419 = ~n_16417 & ~n_16418;
assign n_16420 =  x_636 & ~n_16335;
assign n_16421 =  i_18 &  n_16335;
assign n_16422 = ~n_16420 & ~n_16421;
assign n_16423 =  x_636 & ~n_16422;
assign n_16424 = ~x_636 &  n_16422;
assign n_16425 = ~n_16423 & ~n_16424;
assign n_16426 =  x_635 & ~n_16335;
assign n_16427 =  i_17 &  n_16335;
assign n_16428 = ~n_16426 & ~n_16427;
assign n_16429 =  x_635 & ~n_16428;
assign n_16430 = ~x_635 &  n_16428;
assign n_16431 = ~n_16429 & ~n_16430;
assign n_16432 =  x_634 & ~n_16335;
assign n_16433 =  i_16 &  n_16335;
assign n_16434 = ~n_16432 & ~n_16433;
assign n_16435 =  x_634 & ~n_16434;
assign n_16436 = ~x_634 &  n_16434;
assign n_16437 = ~n_16435 & ~n_16436;
assign n_16438 =  x_633 & ~n_16335;
assign n_16439 =  i_15 &  n_16335;
assign n_16440 = ~n_16438 & ~n_16439;
assign n_16441 =  x_633 & ~n_16440;
assign n_16442 = ~x_633 &  n_16440;
assign n_16443 = ~n_16441 & ~n_16442;
assign n_16444 =  x_632 & ~n_16335;
assign n_16445 =  i_14 &  n_16335;
assign n_16446 = ~n_16444 & ~n_16445;
assign n_16447 =  x_632 & ~n_16446;
assign n_16448 = ~x_632 &  n_16446;
assign n_16449 = ~n_16447 & ~n_16448;
assign n_16450 =  x_631 & ~n_16335;
assign n_16451 =  i_13 &  n_16335;
assign n_16452 = ~n_16450 & ~n_16451;
assign n_16453 =  x_631 & ~n_16452;
assign n_16454 = ~x_631 &  n_16452;
assign n_16455 = ~n_16453 & ~n_16454;
assign n_16456 =  x_630 & ~n_16335;
assign n_16457 =  i_12 &  n_16335;
assign n_16458 = ~n_16456 & ~n_16457;
assign n_16459 =  x_630 & ~n_16458;
assign n_16460 = ~x_630 &  n_16458;
assign n_16461 = ~n_16459 & ~n_16460;
assign n_16462 =  x_629 & ~n_16335;
assign n_16463 =  i_11 &  n_16335;
assign n_16464 = ~n_16462 & ~n_16463;
assign n_16465 =  x_629 & ~n_16464;
assign n_16466 = ~x_629 &  n_16464;
assign n_16467 = ~n_16465 & ~n_16466;
assign n_16468 =  x_628 & ~n_16335;
assign n_16469 =  i_10 &  n_16335;
assign n_16470 = ~n_16468 & ~n_16469;
assign n_16471 =  x_628 & ~n_16470;
assign n_16472 = ~x_628 &  n_16470;
assign n_16473 = ~n_16471 & ~n_16472;
assign n_16474 =  x_627 & ~n_16335;
assign n_16475 =  i_9 &  n_16335;
assign n_16476 = ~n_16474 & ~n_16475;
assign n_16477 =  x_627 & ~n_16476;
assign n_16478 = ~x_627 &  n_16476;
assign n_16479 = ~n_16477 & ~n_16478;
assign n_16480 =  x_626 & ~n_16335;
assign n_16481 =  i_8 &  n_16335;
assign n_16482 = ~n_16480 & ~n_16481;
assign n_16483 =  x_626 & ~n_16482;
assign n_16484 = ~x_626 &  n_16482;
assign n_16485 = ~n_16483 & ~n_16484;
assign n_16486 =  x_625 & ~n_16335;
assign n_16487 =  i_7 &  n_16335;
assign n_16488 = ~n_16486 & ~n_16487;
assign n_16489 =  x_625 & ~n_16488;
assign n_16490 = ~x_625 &  n_16488;
assign n_16491 = ~n_16489 & ~n_16490;
assign n_16492 =  x_624 & ~n_16335;
assign n_16493 =  i_6 &  n_16335;
assign n_16494 = ~n_16492 & ~n_16493;
assign n_16495 =  x_624 & ~n_16494;
assign n_16496 = ~x_624 &  n_16494;
assign n_16497 = ~n_16495 & ~n_16496;
assign n_16498 =  x_623 & ~n_16335;
assign n_16499 =  i_5 &  n_16335;
assign n_16500 = ~n_16498 & ~n_16499;
assign n_16501 =  x_623 & ~n_16500;
assign n_16502 = ~x_623 &  n_16500;
assign n_16503 = ~n_16501 & ~n_16502;
assign n_16504 =  x_622 & ~n_16335;
assign n_16505 =  i_4 &  n_16335;
assign n_16506 = ~n_16504 & ~n_16505;
assign n_16507 =  x_622 & ~n_16506;
assign n_16508 = ~x_622 &  n_16506;
assign n_16509 = ~n_16507 & ~n_16508;
assign n_16510 =  x_621 & ~n_16335;
assign n_16511 =  i_3 &  n_16335;
assign n_16512 = ~n_16510 & ~n_16511;
assign n_16513 =  x_621 & ~n_16512;
assign n_16514 = ~x_621 &  n_16512;
assign n_16515 = ~n_16513 & ~n_16514;
assign n_16516 =  x_620 & ~n_16335;
assign n_16517 =  i_2 &  n_16335;
assign n_16518 = ~n_16516 & ~n_16517;
assign n_16519 =  x_620 & ~n_16518;
assign n_16520 = ~x_620 &  n_16518;
assign n_16521 = ~n_16519 & ~n_16520;
assign n_16522 =  x_619 & ~n_16335;
assign n_16523 =  i_1 &  n_16335;
assign n_16524 = ~n_16522 & ~n_16523;
assign n_16525 =  x_619 & ~n_16524;
assign n_16526 = ~x_619 &  n_16524;
assign n_16527 = ~n_16525 & ~n_16526;
assign n_16528 =  n_980 &  n_1709;
assign n_16529 =  x_618 & ~n_16528;
assign n_16530 =  i_32 &  n_16528;
assign n_16531 = ~n_16529 & ~n_16530;
assign n_16532 =  x_618 & ~n_16531;
assign n_16533 = ~x_618 &  n_16531;
assign n_16534 = ~n_16532 & ~n_16533;
assign n_16535 =  x_617 & ~n_16528;
assign n_16536 =  i_31 &  n_16528;
assign n_16537 = ~n_16535 & ~n_16536;
assign n_16538 =  x_617 & ~n_16537;
assign n_16539 = ~x_617 &  n_16537;
assign n_16540 = ~n_16538 & ~n_16539;
assign n_16541 =  x_616 & ~n_16528;
assign n_16542 =  i_30 &  n_16528;
assign n_16543 = ~n_16541 & ~n_16542;
assign n_16544 =  x_616 & ~n_16543;
assign n_16545 = ~x_616 &  n_16543;
assign n_16546 = ~n_16544 & ~n_16545;
assign n_16547 =  x_615 & ~n_16528;
assign n_16548 =  i_29 &  n_16528;
assign n_16549 = ~n_16547 & ~n_16548;
assign n_16550 =  x_615 & ~n_16549;
assign n_16551 = ~x_615 &  n_16549;
assign n_16552 = ~n_16550 & ~n_16551;
assign n_16553 =  x_614 & ~n_16528;
assign n_16554 =  i_28 &  n_16528;
assign n_16555 = ~n_16553 & ~n_16554;
assign n_16556 =  x_614 & ~n_16555;
assign n_16557 = ~x_614 &  n_16555;
assign n_16558 = ~n_16556 & ~n_16557;
assign n_16559 =  x_613 & ~n_16528;
assign n_16560 =  i_27 &  n_16528;
assign n_16561 = ~n_16559 & ~n_16560;
assign n_16562 =  x_613 & ~n_16561;
assign n_16563 = ~x_613 &  n_16561;
assign n_16564 = ~n_16562 & ~n_16563;
assign n_16565 =  x_612 & ~n_16528;
assign n_16566 =  i_26 &  n_16528;
assign n_16567 = ~n_16565 & ~n_16566;
assign n_16568 =  x_612 & ~n_16567;
assign n_16569 = ~x_612 &  n_16567;
assign n_16570 = ~n_16568 & ~n_16569;
assign n_16571 =  x_611 & ~n_16528;
assign n_16572 =  i_25 &  n_16528;
assign n_16573 = ~n_16571 & ~n_16572;
assign n_16574 =  x_611 & ~n_16573;
assign n_16575 = ~x_611 &  n_16573;
assign n_16576 = ~n_16574 & ~n_16575;
assign n_16577 =  x_610 & ~n_16528;
assign n_16578 =  i_24 &  n_16528;
assign n_16579 = ~n_16577 & ~n_16578;
assign n_16580 =  x_610 & ~n_16579;
assign n_16581 = ~x_610 &  n_16579;
assign n_16582 = ~n_16580 & ~n_16581;
assign n_16583 =  x_609 & ~n_16528;
assign n_16584 =  i_23 &  n_16528;
assign n_16585 = ~n_16583 & ~n_16584;
assign n_16586 =  x_609 & ~n_16585;
assign n_16587 = ~x_609 &  n_16585;
assign n_16588 = ~n_16586 & ~n_16587;
assign n_16589 =  x_608 & ~n_16528;
assign n_16590 =  i_22 &  n_16528;
assign n_16591 = ~n_16589 & ~n_16590;
assign n_16592 =  x_608 & ~n_16591;
assign n_16593 = ~x_608 &  n_16591;
assign n_16594 = ~n_16592 & ~n_16593;
assign n_16595 =  x_607 & ~n_16528;
assign n_16596 =  i_21 &  n_16528;
assign n_16597 = ~n_16595 & ~n_16596;
assign n_16598 =  x_607 & ~n_16597;
assign n_16599 = ~x_607 &  n_16597;
assign n_16600 = ~n_16598 & ~n_16599;
assign n_16601 =  x_606 & ~n_16528;
assign n_16602 =  i_20 &  n_16528;
assign n_16603 = ~n_16601 & ~n_16602;
assign n_16604 =  x_606 & ~n_16603;
assign n_16605 = ~x_606 &  n_16603;
assign n_16606 = ~n_16604 & ~n_16605;
assign n_16607 =  x_605 & ~n_16528;
assign n_16608 =  i_19 &  n_16528;
assign n_16609 = ~n_16607 & ~n_16608;
assign n_16610 =  x_605 & ~n_16609;
assign n_16611 = ~x_605 &  n_16609;
assign n_16612 = ~n_16610 & ~n_16611;
assign n_16613 =  x_604 & ~n_16528;
assign n_16614 =  i_18 &  n_16528;
assign n_16615 = ~n_16613 & ~n_16614;
assign n_16616 =  x_604 & ~n_16615;
assign n_16617 = ~x_604 &  n_16615;
assign n_16618 = ~n_16616 & ~n_16617;
assign n_16619 =  x_603 & ~n_16528;
assign n_16620 =  i_17 &  n_16528;
assign n_16621 = ~n_16619 & ~n_16620;
assign n_16622 =  x_603 & ~n_16621;
assign n_16623 = ~x_603 &  n_16621;
assign n_16624 = ~n_16622 & ~n_16623;
assign n_16625 =  x_602 & ~n_16528;
assign n_16626 =  i_16 &  n_16528;
assign n_16627 = ~n_16625 & ~n_16626;
assign n_16628 =  x_602 & ~n_16627;
assign n_16629 = ~x_602 &  n_16627;
assign n_16630 = ~n_16628 & ~n_16629;
assign n_16631 =  x_601 & ~n_16528;
assign n_16632 =  i_15 &  n_16528;
assign n_16633 = ~n_16631 & ~n_16632;
assign n_16634 =  x_601 & ~n_16633;
assign n_16635 = ~x_601 &  n_16633;
assign n_16636 = ~n_16634 & ~n_16635;
assign n_16637 =  x_600 & ~n_16528;
assign n_16638 =  i_14 &  n_16528;
assign n_16639 = ~n_16637 & ~n_16638;
assign n_16640 =  x_600 & ~n_16639;
assign n_16641 = ~x_600 &  n_16639;
assign n_16642 = ~n_16640 & ~n_16641;
assign n_16643 =  x_599 & ~n_16528;
assign n_16644 =  i_13 &  n_16528;
assign n_16645 = ~n_16643 & ~n_16644;
assign n_16646 =  x_599 & ~n_16645;
assign n_16647 = ~x_599 &  n_16645;
assign n_16648 = ~n_16646 & ~n_16647;
assign n_16649 =  x_598 & ~n_16528;
assign n_16650 =  i_12 &  n_16528;
assign n_16651 = ~n_16649 & ~n_16650;
assign n_16652 =  x_598 & ~n_16651;
assign n_16653 = ~x_598 &  n_16651;
assign n_16654 = ~n_16652 & ~n_16653;
assign n_16655 =  x_597 & ~n_16528;
assign n_16656 =  i_11 &  n_16528;
assign n_16657 = ~n_16655 & ~n_16656;
assign n_16658 =  x_597 & ~n_16657;
assign n_16659 = ~x_597 &  n_16657;
assign n_16660 = ~n_16658 & ~n_16659;
assign n_16661 =  x_596 & ~n_16528;
assign n_16662 =  i_10 &  n_16528;
assign n_16663 = ~n_16661 & ~n_16662;
assign n_16664 =  x_596 & ~n_16663;
assign n_16665 = ~x_596 &  n_16663;
assign n_16666 = ~n_16664 & ~n_16665;
assign n_16667 =  x_595 & ~n_16528;
assign n_16668 =  i_9 &  n_16528;
assign n_16669 = ~n_16667 & ~n_16668;
assign n_16670 =  x_595 & ~n_16669;
assign n_16671 = ~x_595 &  n_16669;
assign n_16672 = ~n_16670 & ~n_16671;
assign n_16673 =  x_594 & ~n_16528;
assign n_16674 =  i_8 &  n_16528;
assign n_16675 = ~n_16673 & ~n_16674;
assign n_16676 =  x_594 & ~n_16675;
assign n_16677 = ~x_594 &  n_16675;
assign n_16678 = ~n_16676 & ~n_16677;
assign n_16679 =  x_593 & ~n_16528;
assign n_16680 =  i_7 &  n_16528;
assign n_16681 = ~n_16679 & ~n_16680;
assign n_16682 =  x_593 & ~n_16681;
assign n_16683 = ~x_593 &  n_16681;
assign n_16684 = ~n_16682 & ~n_16683;
assign n_16685 =  x_592 & ~n_16528;
assign n_16686 =  i_6 &  n_16528;
assign n_16687 = ~n_16685 & ~n_16686;
assign n_16688 =  x_592 & ~n_16687;
assign n_16689 = ~x_592 &  n_16687;
assign n_16690 = ~n_16688 & ~n_16689;
assign n_16691 =  x_591 & ~n_16528;
assign n_16692 =  i_5 &  n_16528;
assign n_16693 = ~n_16691 & ~n_16692;
assign n_16694 =  x_591 & ~n_16693;
assign n_16695 = ~x_591 &  n_16693;
assign n_16696 = ~n_16694 & ~n_16695;
assign n_16697 =  x_590 & ~n_16528;
assign n_16698 =  i_4 &  n_16528;
assign n_16699 = ~n_16697 & ~n_16698;
assign n_16700 =  x_590 & ~n_16699;
assign n_16701 = ~x_590 &  n_16699;
assign n_16702 = ~n_16700 & ~n_16701;
assign n_16703 =  x_589 & ~n_16528;
assign n_16704 =  i_3 &  n_16528;
assign n_16705 = ~n_16703 & ~n_16704;
assign n_16706 =  x_589 & ~n_16705;
assign n_16707 = ~x_589 &  n_16705;
assign n_16708 = ~n_16706 & ~n_16707;
assign n_16709 =  x_588 & ~n_16528;
assign n_16710 =  i_2 &  n_16528;
assign n_16711 = ~n_16709 & ~n_16710;
assign n_16712 =  x_588 & ~n_16711;
assign n_16713 = ~x_588 &  n_16711;
assign n_16714 = ~n_16712 & ~n_16713;
assign n_16715 =  x_587 & ~n_16528;
assign n_16716 =  i_1 &  n_16528;
assign n_16717 = ~n_16715 & ~n_16716;
assign n_16718 =  x_587 & ~n_16717;
assign n_16719 = ~x_587 &  n_16717;
assign n_16720 = ~n_16718 & ~n_16719;
assign n_16721 =  n_6532 &  n_980;
assign n_16722 =  x_586 & ~n_16721;
assign n_16723 =  i_32 &  n_16721;
assign n_16724 = ~n_16722 & ~n_16723;
assign n_16725 =  x_586 & ~n_16724;
assign n_16726 = ~x_586 &  n_16724;
assign n_16727 = ~n_16725 & ~n_16726;
assign n_16728 =  x_585 & ~n_16721;
assign n_16729 =  i_31 &  n_16721;
assign n_16730 = ~n_16728 & ~n_16729;
assign n_16731 =  x_585 & ~n_16730;
assign n_16732 = ~x_585 &  n_16730;
assign n_16733 = ~n_16731 & ~n_16732;
assign n_16734 =  x_584 & ~n_16721;
assign n_16735 =  i_30 &  n_16721;
assign n_16736 = ~n_16734 & ~n_16735;
assign n_16737 =  x_584 & ~n_16736;
assign n_16738 = ~x_584 &  n_16736;
assign n_16739 = ~n_16737 & ~n_16738;
assign n_16740 =  x_583 & ~n_16721;
assign n_16741 =  i_29 &  n_16721;
assign n_16742 = ~n_16740 & ~n_16741;
assign n_16743 =  x_583 & ~n_16742;
assign n_16744 = ~x_583 &  n_16742;
assign n_16745 = ~n_16743 & ~n_16744;
assign n_16746 =  x_582 & ~n_16721;
assign n_16747 =  i_28 &  n_16721;
assign n_16748 = ~n_16746 & ~n_16747;
assign n_16749 =  x_582 & ~n_16748;
assign n_16750 = ~x_582 &  n_16748;
assign n_16751 = ~n_16749 & ~n_16750;
assign n_16752 =  x_581 & ~n_16721;
assign n_16753 =  i_27 &  n_16721;
assign n_16754 = ~n_16752 & ~n_16753;
assign n_16755 =  x_581 & ~n_16754;
assign n_16756 = ~x_581 &  n_16754;
assign n_16757 = ~n_16755 & ~n_16756;
assign n_16758 =  x_580 & ~n_16721;
assign n_16759 =  i_26 &  n_16721;
assign n_16760 = ~n_16758 & ~n_16759;
assign n_16761 =  x_580 & ~n_16760;
assign n_16762 = ~x_580 &  n_16760;
assign n_16763 = ~n_16761 & ~n_16762;
assign n_16764 =  x_579 & ~n_16721;
assign n_16765 =  i_25 &  n_16721;
assign n_16766 = ~n_16764 & ~n_16765;
assign n_16767 =  x_579 & ~n_16766;
assign n_16768 = ~x_579 &  n_16766;
assign n_16769 = ~n_16767 & ~n_16768;
assign n_16770 =  x_578 & ~n_16721;
assign n_16771 =  i_24 &  n_16721;
assign n_16772 = ~n_16770 & ~n_16771;
assign n_16773 =  x_578 & ~n_16772;
assign n_16774 = ~x_578 &  n_16772;
assign n_16775 = ~n_16773 & ~n_16774;
assign n_16776 =  x_577 & ~n_16721;
assign n_16777 =  i_23 &  n_16721;
assign n_16778 = ~n_16776 & ~n_16777;
assign n_16779 =  x_577 & ~n_16778;
assign n_16780 = ~x_577 &  n_16778;
assign n_16781 = ~n_16779 & ~n_16780;
assign n_16782 =  x_576 & ~n_16721;
assign n_16783 =  i_22 &  n_16721;
assign n_16784 = ~n_16782 & ~n_16783;
assign n_16785 =  x_576 & ~n_16784;
assign n_16786 = ~x_576 &  n_16784;
assign n_16787 = ~n_16785 & ~n_16786;
assign n_16788 =  x_575 & ~n_16721;
assign n_16789 =  i_21 &  n_16721;
assign n_16790 = ~n_16788 & ~n_16789;
assign n_16791 =  x_575 & ~n_16790;
assign n_16792 = ~x_575 &  n_16790;
assign n_16793 = ~n_16791 & ~n_16792;
assign n_16794 =  x_574 & ~n_16721;
assign n_16795 =  i_20 &  n_16721;
assign n_16796 = ~n_16794 & ~n_16795;
assign n_16797 =  x_574 & ~n_16796;
assign n_16798 = ~x_574 &  n_16796;
assign n_16799 = ~n_16797 & ~n_16798;
assign n_16800 =  x_573 & ~n_16721;
assign n_16801 =  i_19 &  n_16721;
assign n_16802 = ~n_16800 & ~n_16801;
assign n_16803 =  x_573 & ~n_16802;
assign n_16804 = ~x_573 &  n_16802;
assign n_16805 = ~n_16803 & ~n_16804;
assign n_16806 =  x_572 & ~n_16721;
assign n_16807 =  i_18 &  n_16721;
assign n_16808 = ~n_16806 & ~n_16807;
assign n_16809 =  x_572 & ~n_16808;
assign n_16810 = ~x_572 &  n_16808;
assign n_16811 = ~n_16809 & ~n_16810;
assign n_16812 =  x_571 & ~n_16721;
assign n_16813 =  i_17 &  n_16721;
assign n_16814 = ~n_16812 & ~n_16813;
assign n_16815 =  x_571 & ~n_16814;
assign n_16816 = ~x_571 &  n_16814;
assign n_16817 = ~n_16815 & ~n_16816;
assign n_16818 =  x_570 & ~n_16721;
assign n_16819 =  i_16 &  n_16721;
assign n_16820 = ~n_16818 & ~n_16819;
assign n_16821 =  x_570 & ~n_16820;
assign n_16822 = ~x_570 &  n_16820;
assign n_16823 = ~n_16821 & ~n_16822;
assign n_16824 =  x_569 & ~n_16721;
assign n_16825 =  i_15 &  n_16721;
assign n_16826 = ~n_16824 & ~n_16825;
assign n_16827 =  x_569 & ~n_16826;
assign n_16828 = ~x_569 &  n_16826;
assign n_16829 = ~n_16827 & ~n_16828;
assign n_16830 =  x_568 & ~n_16721;
assign n_16831 =  i_14 &  n_16721;
assign n_16832 = ~n_16830 & ~n_16831;
assign n_16833 =  x_568 & ~n_16832;
assign n_16834 = ~x_568 &  n_16832;
assign n_16835 = ~n_16833 & ~n_16834;
assign n_16836 =  x_567 & ~n_16721;
assign n_16837 =  i_13 &  n_16721;
assign n_16838 = ~n_16836 & ~n_16837;
assign n_16839 =  x_567 & ~n_16838;
assign n_16840 = ~x_567 &  n_16838;
assign n_16841 = ~n_16839 & ~n_16840;
assign n_16842 =  x_566 & ~n_16721;
assign n_16843 =  i_12 &  n_16721;
assign n_16844 = ~n_16842 & ~n_16843;
assign n_16845 =  x_566 & ~n_16844;
assign n_16846 = ~x_566 &  n_16844;
assign n_16847 = ~n_16845 & ~n_16846;
assign n_16848 =  x_565 & ~n_16721;
assign n_16849 =  i_11 &  n_16721;
assign n_16850 = ~n_16848 & ~n_16849;
assign n_16851 =  x_565 & ~n_16850;
assign n_16852 = ~x_565 &  n_16850;
assign n_16853 = ~n_16851 & ~n_16852;
assign n_16854 =  x_564 & ~n_16721;
assign n_16855 =  i_10 &  n_16721;
assign n_16856 = ~n_16854 & ~n_16855;
assign n_16857 =  x_564 & ~n_16856;
assign n_16858 = ~x_564 &  n_16856;
assign n_16859 = ~n_16857 & ~n_16858;
assign n_16860 =  x_563 & ~n_16721;
assign n_16861 =  i_9 &  n_16721;
assign n_16862 = ~n_16860 & ~n_16861;
assign n_16863 =  x_563 & ~n_16862;
assign n_16864 = ~x_563 &  n_16862;
assign n_16865 = ~n_16863 & ~n_16864;
assign n_16866 =  x_562 & ~n_16721;
assign n_16867 =  i_8 &  n_16721;
assign n_16868 = ~n_16866 & ~n_16867;
assign n_16869 =  x_562 & ~n_16868;
assign n_16870 = ~x_562 &  n_16868;
assign n_16871 = ~n_16869 & ~n_16870;
assign n_16872 =  x_561 & ~n_16721;
assign n_16873 =  i_7 &  n_16721;
assign n_16874 = ~n_16872 & ~n_16873;
assign n_16875 =  x_561 & ~n_16874;
assign n_16876 = ~x_561 &  n_16874;
assign n_16877 = ~n_16875 & ~n_16876;
assign n_16878 =  x_560 & ~n_16721;
assign n_16879 =  i_6 &  n_16721;
assign n_16880 = ~n_16878 & ~n_16879;
assign n_16881 =  x_560 & ~n_16880;
assign n_16882 = ~x_560 &  n_16880;
assign n_16883 = ~n_16881 & ~n_16882;
assign n_16884 =  x_559 & ~n_16721;
assign n_16885 =  i_5 &  n_16721;
assign n_16886 = ~n_16884 & ~n_16885;
assign n_16887 =  x_559 & ~n_16886;
assign n_16888 = ~x_559 &  n_16886;
assign n_16889 = ~n_16887 & ~n_16888;
assign n_16890 =  x_558 & ~n_16721;
assign n_16891 =  i_4 &  n_16721;
assign n_16892 = ~n_16890 & ~n_16891;
assign n_16893 =  x_558 & ~n_16892;
assign n_16894 = ~x_558 &  n_16892;
assign n_16895 = ~n_16893 & ~n_16894;
assign n_16896 =  x_557 & ~n_16721;
assign n_16897 =  i_3 &  n_16721;
assign n_16898 = ~n_16896 & ~n_16897;
assign n_16899 =  x_557 & ~n_16898;
assign n_16900 = ~x_557 &  n_16898;
assign n_16901 = ~n_16899 & ~n_16900;
assign n_16902 =  x_556 & ~n_16721;
assign n_16903 =  i_2 &  n_16721;
assign n_16904 = ~n_16902 & ~n_16903;
assign n_16905 =  x_556 & ~n_16904;
assign n_16906 = ~x_556 &  n_16904;
assign n_16907 = ~n_16905 & ~n_16906;
assign n_16908 =  x_555 & ~n_16721;
assign n_16909 =  i_1 &  n_16721;
assign n_16910 = ~n_16908 & ~n_16909;
assign n_16911 =  x_555 & ~n_16910;
assign n_16912 = ~x_555 &  n_16910;
assign n_16913 = ~n_16911 & ~n_16912;
assign n_16914 =  x_39 &  n_12226;
assign n_16915 = ~n_2499 & ~n_4251;
assign n_16916 = ~n_16914 &  n_16915;
assign n_16917 =  n_12614 & ~n_16916;
assign n_16918 =  x_554 & ~n_16917;
assign n_16919 =  n_2499 &  n_12614;
assign n_16920 = ~x_39 &  n_16919;
assign n_16921 =  x_74 &  x_1962;
assign n_16922 = ~x_74 & ~x_1962;
assign n_16923 = ~n_16921 & ~n_16922;
assign n_16924 =  n_16920 &  n_16923;
assign n_16925 =  n_8254 &  n_12226;
assign n_16926 =  x_1034 &  n_16925;
assign n_16927 =  n_12614 &  n_4251;
assign n_16928 =  x_298 &  x_1674;
assign n_16929 = ~x_298 & ~x_1674;
assign n_16930 = ~n_16928 & ~n_16929;
assign n_16931 =  n_16927 &  n_16930;
assign n_16932 =  n_8254 &  n_2499;
assign n_16933 =  x_2570 &  x_2634;
assign n_16934 = ~x_2570 & ~x_2634;
assign n_16935 = ~n_16933 & ~n_16934;
assign n_16936 =  n_16932 &  n_16935;
assign n_16937 = ~n_16931 & ~n_16936;
assign n_16938 = ~n_16926 &  n_16937;
assign n_16939 = ~n_16924 &  n_16938;
assign n_16940 = ~n_16918 &  n_16939;
assign n_16941 =  x_554 & ~n_16940;
assign n_16942 = ~x_554 &  n_16940;
assign n_16943 = ~n_16941 & ~n_16942;
assign n_16944 =  x_553 & ~n_16917;
assign n_16945 = ~x_2633 & ~x_2634;
assign n_16946 =  x_2633 &  x_2634;
assign n_16947 = ~n_16945 & ~n_16946;
assign n_16948 =  x_2569 &  n_16947;
assign n_16949 = ~x_2569 & ~n_16947;
assign n_16950 = ~n_16948 & ~n_16949;
assign n_16951 = ~n_16933 & ~n_16950;
assign n_16952 =  n_16933 &  n_16950;
assign n_16953 =  n_16932 & ~n_16952;
assign n_16954 = ~n_16951 &  n_16953;
assign n_16955 = ~x_1033 & ~x_1034;
assign n_16956 =  x_1033 &  x_1034;
assign n_16957 = ~n_16955 & ~n_16956;
assign n_16958 =  n_16925 &  n_16957;
assign n_16959 = ~n_16954 & ~n_16958;
assign n_16960 = ~x_73 & ~x_74;
assign n_16961 =  x_73 &  x_74;
assign n_16962 = ~n_16960 & ~n_16961;
assign n_16963 =  x_1961 &  n_16962;
assign n_16964 = ~x_1961 & ~n_16962;
assign n_16965 = ~n_16963 & ~n_16964;
assign n_16966 =  n_16921 &  n_16965;
assign n_16967 = ~n_16921 & ~n_16965;
assign n_16968 = ~n_16966 & ~n_16967;
assign n_16969 =  n_16920 &  n_16968;
assign n_16970 = ~x_1673 & ~x_1674;
assign n_16971 =  x_1673 &  x_1674;
assign n_16972 = ~n_16970 & ~n_16971;
assign n_16973 =  x_297 &  n_16972;
assign n_16974 = ~x_297 & ~n_16972;
assign n_16975 = ~n_16973 & ~n_16974;
assign n_16976 = ~n_16928 & ~n_16975;
assign n_16977 =  n_16928 &  n_16975;
assign n_16978 =  n_16927 & ~n_16977;
assign n_16979 = ~n_16976 &  n_16978;
assign n_16980 = ~n_16969 & ~n_16979;
assign n_16981 =  n_16959 &  n_16980;
assign n_16982 = ~n_16944 &  n_16981;
assign n_16983 =  x_553 & ~n_16982;
assign n_16984 = ~x_553 &  n_16982;
assign n_16985 = ~n_16983 & ~n_16984;
assign n_16986 =  x_552 & ~n_16917;
assign n_16987 = ~x_1032 &  n_16955;
assign n_16988 =  x_1032 & ~n_16955;
assign n_16989 = ~n_16987 & ~n_16988;
assign n_16990 =  n_16925 &  n_16989;
assign n_16991 = ~n_16986 & ~n_16990;
assign n_16992 = ~x_2632 &  n_16945;
assign n_16993 =  x_2632 & ~n_16945;
assign n_16994 = ~n_16992 & ~n_16993;
assign n_16995 = ~x_2569 &  x_2633;
assign n_16996 =  n_16933 & ~n_16995;
assign n_16997 = ~n_16996 & ~n_16948;
assign n_16998 =  n_16994 & ~n_16997;
assign n_16999 = ~n_16994 &  n_16997;
assign n_17000 = ~n_16998 & ~n_16999;
assign n_17001 = ~x_2568 & ~n_17000;
assign n_17002 =  x_2568 & ~n_16999;
assign n_17003 = ~n_16998 &  n_17002;
assign n_17004 =  n_16932 & ~n_17003;
assign n_17005 = ~n_17001 &  n_17004;
assign n_17006 = ~x_1672 &  n_16970;
assign n_17007 =  x_1672 & ~n_16970;
assign n_17008 = ~n_17006 & ~n_17007;
assign n_17009 = ~x_297 &  x_1673;
assign n_17010 =  n_16928 & ~n_17009;
assign n_17011 = ~n_17010 & ~n_16973;
assign n_17012 =  n_17008 & ~n_17011;
assign n_17013 = ~n_17008 &  n_17011;
assign n_17014 = ~n_17012 & ~n_17013;
assign n_17015 = ~x_296 & ~n_17014;
assign n_17016 =  x_296 & ~n_17013;
assign n_17017 = ~n_17012 &  n_17016;
assign n_17018 =  n_16927 & ~n_17017;
assign n_17019 = ~n_17015 &  n_17018;
assign n_17020 = ~x_72 &  n_16960;
assign n_17021 =  x_72 & ~n_16960;
assign n_17022 = ~n_17020 & ~n_17021;
assign n_17023 =  x_73 & ~x_1961;
assign n_17024 =  n_16921 & ~n_17023;
assign n_17025 = ~n_17024 & ~n_16963;
assign n_17026 =  n_17022 & ~n_17025;
assign n_17027 = ~n_17022 &  n_17025;
assign n_17028 = ~n_17026 & ~n_17027;
assign n_17029 = ~x_1960 & ~n_17028;
assign n_17030 =  x_1960 & ~n_17027;
assign n_17031 = ~n_17026 &  n_17030;
assign n_17032 =  n_16920 & ~n_17031;
assign n_17033 = ~n_17029 &  n_17032;
assign n_17034 = ~n_17019 & ~n_17033;
assign n_17035 = ~n_17005 &  n_17034;
assign n_17036 =  n_16991 &  n_17035;
assign n_17037 =  x_552 & ~n_17036;
assign n_17038 = ~x_552 &  n_17036;
assign n_17039 = ~n_17037 & ~n_17038;
assign n_17040 = ~x_1671 &  n_17006;
assign n_17041 =  x_1671 & ~n_17006;
assign n_17042 = ~n_17040 & ~n_17041;
assign n_17043 = ~n_17012 & ~n_17016;
assign n_17044 =  n_17042 & ~n_17043;
assign n_17045 = ~n_17042 &  n_17043;
assign n_17046 = ~n_17044 & ~n_17045;
assign n_17047 = ~x_295 & ~n_17046;
assign n_17048 =  x_295 & ~n_17045;
assign n_17049 = ~n_17044 &  n_17048;
assign n_17050 =  n_16927 & ~n_17049;
assign n_17051 = ~n_17047 &  n_17050;
assign n_17052 =  x_551 & ~n_16917;
assign n_17053 = ~x_1031 &  n_16987;
assign n_17054 =  x_1031 & ~n_16987;
assign n_17055 = ~n_17053 & ~n_17054;
assign n_17056 =  n_16925 &  n_17055;
assign n_17057 = ~n_17052 & ~n_17056;
assign n_17058 = ~n_17051 &  n_17057;
assign n_17059 = ~x_71 &  n_17020;
assign n_17060 =  x_71 & ~n_17020;
assign n_17061 = ~n_17059 & ~n_17060;
assign n_17062 = ~n_17026 & ~n_17030;
assign n_17063 =  n_17061 & ~n_17062;
assign n_17064 = ~n_17061 &  n_17062;
assign n_17065 = ~n_17063 & ~n_17064;
assign n_17066 = ~x_1959 & ~n_17065;
assign n_17067 =  x_1959 & ~n_17064;
assign n_17068 = ~n_17063 &  n_17067;
assign n_17069 =  n_16920 & ~n_17068;
assign n_17070 = ~n_17066 &  n_17069;
assign n_17071 = ~x_2631 &  n_16992;
assign n_17072 =  x_2631 & ~n_16992;
assign n_17073 = ~n_17071 & ~n_17072;
assign n_17074 = ~n_16998 & ~n_17002;
assign n_17075 =  n_17073 & ~n_17074;
assign n_17076 = ~n_17073 &  n_17074;
assign n_17077 = ~n_17075 & ~n_17076;
assign n_17078 = ~x_2567 & ~n_17077;
assign n_17079 =  x_2567 & ~n_17076;
assign n_17080 = ~n_17075 &  n_17079;
assign n_17081 =  n_16932 & ~n_17080;
assign n_17082 = ~n_17078 &  n_17081;
assign n_17083 = ~n_17070 & ~n_17082;
assign n_17084 =  n_17058 &  n_17083;
assign n_17085 =  x_551 & ~n_17084;
assign n_17086 = ~x_551 &  n_17084;
assign n_17087 = ~n_17085 & ~n_17086;
assign n_17088 = ~x_1670 &  n_17040;
assign n_17089 =  x_1670 & ~n_17040;
assign n_17090 = ~n_17088 & ~n_17089;
assign n_17091 = ~n_17044 & ~n_17048;
assign n_17092 =  n_17090 & ~n_17091;
assign n_17093 = ~n_17090 &  n_17091;
assign n_17094 = ~n_17092 & ~n_17093;
assign n_17095 = ~x_294 & ~n_17094;
assign n_17096 =  x_294 & ~n_17093;
assign n_17097 = ~n_17092 &  n_17096;
assign n_17098 =  n_16927 & ~n_17097;
assign n_17099 = ~n_17095 &  n_17098;
assign n_17100 =  x_550 & ~n_16917;
assign n_17101 = ~x_1030 &  n_17053;
assign n_17102 =  x_1030 & ~n_17053;
assign n_17103 = ~n_17101 & ~n_17102;
assign n_17104 =  n_16925 &  n_17103;
assign n_17105 = ~n_17100 & ~n_17104;
assign n_17106 = ~n_17099 &  n_17105;
assign n_17107 = ~x_70 &  n_17059;
assign n_17108 =  x_70 & ~n_17059;
assign n_17109 = ~n_17107 & ~n_17108;
assign n_17110 = ~n_17063 & ~n_17067;
assign n_17111 =  n_17109 & ~n_17110;
assign n_17112 = ~n_17109 &  n_17110;
assign n_17113 = ~n_17111 & ~n_17112;
assign n_17114 = ~x_1958 & ~n_17113;
assign n_17115 =  x_1958 & ~n_17112;
assign n_17116 = ~n_17111 &  n_17115;
assign n_17117 =  n_16920 & ~n_17116;
assign n_17118 = ~n_17114 &  n_17117;
assign n_17119 = ~x_2630 &  n_17071;
assign n_17120 =  x_2630 & ~n_17071;
assign n_17121 = ~n_17119 & ~n_17120;
assign n_17122 = ~n_17075 & ~n_17079;
assign n_17123 =  n_17121 & ~n_17122;
assign n_17124 = ~n_17121 &  n_17122;
assign n_17125 = ~n_17123 & ~n_17124;
assign n_17126 = ~x_2566 & ~n_17125;
assign n_17127 =  x_2566 & ~n_17124;
assign n_17128 = ~n_17123 &  n_17127;
assign n_17129 =  n_16932 & ~n_17128;
assign n_17130 = ~n_17126 &  n_17129;
assign n_17131 = ~n_17118 & ~n_17130;
assign n_17132 =  n_17106 &  n_17131;
assign n_17133 =  x_550 & ~n_17132;
assign n_17134 = ~x_550 &  n_17132;
assign n_17135 = ~n_17133 & ~n_17134;
assign n_17136 = ~x_1669 &  n_17088;
assign n_17137 =  x_1669 & ~n_17088;
assign n_17138 = ~n_17136 & ~n_17137;
assign n_17139 = ~n_17092 & ~n_17096;
assign n_17140 =  n_17138 & ~n_17139;
assign n_17141 = ~n_17138 &  n_17139;
assign n_17142 = ~n_17140 & ~n_17141;
assign n_17143 = ~x_293 & ~n_17142;
assign n_17144 =  x_293 & ~n_17141;
assign n_17145 = ~n_17140 &  n_17144;
assign n_17146 =  n_16927 & ~n_17145;
assign n_17147 = ~n_17143 &  n_17146;
assign n_17148 =  x_549 & ~n_16917;
assign n_17149 = ~x_1029 &  n_17101;
assign n_17150 =  x_1029 & ~n_17101;
assign n_17151 = ~n_17149 & ~n_17150;
assign n_17152 =  n_16925 &  n_17151;
assign n_17153 = ~n_17148 & ~n_17152;
assign n_17154 = ~n_17147 &  n_17153;
assign n_17155 = ~x_69 &  n_17107;
assign n_17156 =  x_69 & ~n_17107;
assign n_17157 = ~n_17155 & ~n_17156;
assign n_17158 = ~n_17111 & ~n_17115;
assign n_17159 =  n_17157 & ~n_17158;
assign n_17160 = ~n_17157 &  n_17158;
assign n_17161 = ~n_17159 & ~n_17160;
assign n_17162 = ~x_1957 & ~n_17161;
assign n_17163 =  x_1957 & ~n_17160;
assign n_17164 = ~n_17159 &  n_17163;
assign n_17165 =  n_16920 & ~n_17164;
assign n_17166 = ~n_17162 &  n_17165;
assign n_17167 = ~x_2629 &  n_17119;
assign n_17168 =  x_2629 & ~n_17119;
assign n_17169 = ~n_17167 & ~n_17168;
assign n_17170 = ~n_17123 & ~n_17127;
assign n_17171 =  n_17169 & ~n_17170;
assign n_17172 = ~n_17169 &  n_17170;
assign n_17173 = ~n_17171 & ~n_17172;
assign n_17174 = ~x_2565 & ~n_17173;
assign n_17175 =  x_2565 & ~n_17172;
assign n_17176 = ~n_17171 &  n_17175;
assign n_17177 =  n_16932 & ~n_17176;
assign n_17178 = ~n_17174 &  n_17177;
assign n_17179 = ~n_17166 & ~n_17178;
assign n_17180 =  n_17154 &  n_17179;
assign n_17181 =  x_549 & ~n_17180;
assign n_17182 = ~x_549 &  n_17180;
assign n_17183 = ~n_17181 & ~n_17182;
assign n_17184 = ~x_1668 &  n_17136;
assign n_17185 =  x_1668 & ~n_17136;
assign n_17186 = ~n_17184 & ~n_17185;
assign n_17187 = ~n_17140 & ~n_17144;
assign n_17188 =  n_17186 & ~n_17187;
assign n_17189 = ~n_17186 &  n_17187;
assign n_17190 = ~n_17188 & ~n_17189;
assign n_17191 = ~x_292 & ~n_17190;
assign n_17192 =  x_292 & ~n_17189;
assign n_17193 = ~n_17188 &  n_17192;
assign n_17194 =  n_16927 & ~n_17193;
assign n_17195 = ~n_17191 &  n_17194;
assign n_17196 =  x_548 & ~n_16917;
assign n_17197 =  x_1028 & ~n_17149;
assign n_17198 = ~x_1028 &  n_17149;
assign n_17199 =  n_16925 & ~n_17198;
assign n_17200 = ~n_17197 &  n_17199;
assign n_17201 = ~n_17196 & ~n_17200;
assign n_17202 = ~n_17195 &  n_17201;
assign n_17203 = ~x_68 &  n_17155;
assign n_17204 =  x_68 & ~n_17155;
assign n_17205 = ~n_17203 & ~n_17204;
assign n_17206 = ~n_17159 & ~n_17163;
assign n_17207 =  n_17205 & ~n_17206;
assign n_17208 = ~n_17205 &  n_17206;
assign n_17209 = ~n_17207 & ~n_17208;
assign n_17210 = ~x_1956 & ~n_17209;
assign n_17211 =  x_1956 & ~n_17208;
assign n_17212 = ~n_17207 &  n_17211;
assign n_17213 =  n_16920 & ~n_17212;
assign n_17214 = ~n_17210 &  n_17213;
assign n_17215 = ~x_2628 &  n_17167;
assign n_17216 =  x_2628 & ~n_17167;
assign n_17217 = ~n_17215 & ~n_17216;
assign n_17218 = ~n_17171 & ~n_17175;
assign n_17219 =  n_17217 & ~n_17218;
assign n_17220 = ~n_17217 &  n_17218;
assign n_17221 = ~n_17219 & ~n_17220;
assign n_17222 = ~x_2564 & ~n_17221;
assign n_17223 =  x_2564 & ~n_17220;
assign n_17224 = ~n_17219 &  n_17223;
assign n_17225 =  n_16932 & ~n_17224;
assign n_17226 = ~n_17222 &  n_17225;
assign n_17227 = ~n_17214 & ~n_17226;
assign n_17228 =  n_17202 &  n_17227;
assign n_17229 =  x_548 & ~n_17228;
assign n_17230 = ~x_548 &  n_17228;
assign n_17231 = ~n_17229 & ~n_17230;
assign n_17232 = ~x_1667 &  n_17184;
assign n_17233 =  x_1667 & ~n_17184;
assign n_17234 = ~n_17232 & ~n_17233;
assign n_17235 = ~n_17188 & ~n_17192;
assign n_17236 =  n_17234 & ~n_17235;
assign n_17237 = ~n_17234 &  n_17235;
assign n_17238 = ~n_17236 & ~n_17237;
assign n_17239 = ~x_291 & ~n_17238;
assign n_17240 =  x_291 & ~n_17237;
assign n_17241 = ~n_17236 &  n_17240;
assign n_17242 =  n_16927 & ~n_17241;
assign n_17243 = ~n_17239 &  n_17242;
assign n_17244 =  x_547 & ~n_16917;
assign n_17245 =  x_1027 & ~n_17198;
assign n_17246 = ~x_1027 &  n_17198;
assign n_17247 =  n_16925 & ~n_17246;
assign n_17248 = ~n_17245 &  n_17247;
assign n_17249 = ~n_17244 & ~n_17248;
assign n_17250 = ~n_17243 &  n_17249;
assign n_17251 = ~x_67 &  n_17203;
assign n_17252 =  x_67 & ~n_17203;
assign n_17253 = ~n_17251 & ~n_17252;
assign n_17254 = ~n_17207 & ~n_17211;
assign n_17255 =  n_17253 & ~n_17254;
assign n_17256 = ~n_17253 &  n_17254;
assign n_17257 = ~n_17255 & ~n_17256;
assign n_17258 = ~x_1955 & ~n_17257;
assign n_17259 =  x_1955 & ~n_17256;
assign n_17260 = ~n_17255 &  n_17259;
assign n_17261 =  n_16920 & ~n_17260;
assign n_17262 = ~n_17258 &  n_17261;
assign n_17263 = ~x_2627 &  n_17215;
assign n_17264 =  x_2627 & ~n_17215;
assign n_17265 = ~n_17263 & ~n_17264;
assign n_17266 = ~n_17219 & ~n_17223;
assign n_17267 =  n_17265 & ~n_17266;
assign n_17268 = ~n_17265 &  n_17266;
assign n_17269 = ~n_17267 & ~n_17268;
assign n_17270 = ~x_2563 & ~n_17269;
assign n_17271 =  x_2563 & ~n_17268;
assign n_17272 = ~n_17267 &  n_17271;
assign n_17273 =  n_16932 & ~n_17272;
assign n_17274 = ~n_17270 &  n_17273;
assign n_17275 = ~n_17262 & ~n_17274;
assign n_17276 =  n_17250 &  n_17275;
assign n_17277 =  x_547 & ~n_17276;
assign n_17278 = ~x_547 &  n_17276;
assign n_17279 = ~n_17277 & ~n_17278;
assign n_17280 = ~x_1666 &  n_17232;
assign n_17281 =  x_1666 & ~n_17232;
assign n_17282 = ~n_17280 & ~n_17281;
assign n_17283 = ~n_17236 & ~n_17240;
assign n_17284 =  n_17282 & ~n_17283;
assign n_17285 = ~n_17282 &  n_17283;
assign n_17286 = ~n_17284 & ~n_17285;
assign n_17287 = ~x_290 & ~n_17286;
assign n_17288 =  x_290 & ~n_17285;
assign n_17289 = ~n_17284 &  n_17288;
assign n_17290 =  n_16927 & ~n_17289;
assign n_17291 = ~n_17287 &  n_17290;
assign n_17292 =  x_546 & ~n_16917;
assign n_17293 =  x_1026 & ~n_17246;
assign n_17294 = ~x_1026 &  n_17246;
assign n_17295 =  n_16925 & ~n_17294;
assign n_17296 = ~n_17293 &  n_17295;
assign n_17297 = ~n_17292 & ~n_17296;
assign n_17298 = ~n_17291 &  n_17297;
assign n_17299 = ~x_66 &  n_17251;
assign n_17300 =  x_66 & ~n_17251;
assign n_17301 = ~n_17299 & ~n_17300;
assign n_17302 = ~n_17255 & ~n_17259;
assign n_17303 =  n_17301 & ~n_17302;
assign n_17304 = ~n_17301 &  n_17302;
assign n_17305 = ~n_17303 & ~n_17304;
assign n_17306 = ~x_1954 & ~n_17305;
assign n_17307 =  x_1954 & ~n_17304;
assign n_17308 = ~n_17303 &  n_17307;
assign n_17309 =  n_16920 & ~n_17308;
assign n_17310 = ~n_17306 &  n_17309;
assign n_17311 = ~x_2626 &  n_17263;
assign n_17312 =  x_2626 & ~n_17263;
assign n_17313 = ~n_17311 & ~n_17312;
assign n_17314 = ~n_17267 & ~n_17271;
assign n_17315 =  n_17313 & ~n_17314;
assign n_17316 = ~n_17313 &  n_17314;
assign n_17317 = ~n_17315 & ~n_17316;
assign n_17318 = ~x_2562 & ~n_17317;
assign n_17319 =  x_2562 & ~n_17316;
assign n_17320 = ~n_17315 &  n_17319;
assign n_17321 =  n_16932 & ~n_17320;
assign n_17322 = ~n_17318 &  n_17321;
assign n_17323 = ~n_17310 & ~n_17322;
assign n_17324 =  n_17298 &  n_17323;
assign n_17325 =  x_546 & ~n_17324;
assign n_17326 = ~x_546 &  n_17324;
assign n_17327 = ~n_17325 & ~n_17326;
assign n_17328 = ~x_1665 &  n_17280;
assign n_17329 =  x_1665 & ~n_17280;
assign n_17330 = ~n_17328 & ~n_17329;
assign n_17331 = ~n_17284 & ~n_17288;
assign n_17332 =  n_17330 & ~n_17331;
assign n_17333 = ~n_17330 &  n_17331;
assign n_17334 = ~n_17332 & ~n_17333;
assign n_17335 = ~x_289 & ~n_17334;
assign n_17336 =  x_289 & ~n_17333;
assign n_17337 = ~n_17332 &  n_17336;
assign n_17338 =  n_16927 & ~n_17337;
assign n_17339 = ~n_17335 &  n_17338;
assign n_17340 =  x_545 & ~n_16917;
assign n_17341 =  x_1025 & ~n_17294;
assign n_17342 = ~x_1025 &  n_17294;
assign n_17343 =  n_16925 & ~n_17342;
assign n_17344 = ~n_17341 &  n_17343;
assign n_17345 = ~n_17340 & ~n_17344;
assign n_17346 = ~n_17339 &  n_17345;
assign n_17347 = ~x_65 &  n_17299;
assign n_17348 =  x_65 & ~n_17299;
assign n_17349 = ~n_17347 & ~n_17348;
assign n_17350 = ~n_17303 & ~n_17307;
assign n_17351 =  n_17349 & ~n_17350;
assign n_17352 = ~n_17349 &  n_17350;
assign n_17353 = ~n_17351 & ~n_17352;
assign n_17354 = ~x_1953 & ~n_17353;
assign n_17355 =  x_1953 & ~n_17352;
assign n_17356 = ~n_17351 &  n_17355;
assign n_17357 =  n_16920 & ~n_17356;
assign n_17358 = ~n_17354 &  n_17357;
assign n_17359 = ~x_2625 &  n_17311;
assign n_17360 =  x_2625 & ~n_17311;
assign n_17361 = ~n_17359 & ~n_17360;
assign n_17362 = ~n_17315 & ~n_17319;
assign n_17363 =  n_17361 & ~n_17362;
assign n_17364 = ~n_17361 &  n_17362;
assign n_17365 = ~n_17363 & ~n_17364;
assign n_17366 = ~x_2561 & ~n_17365;
assign n_17367 =  x_2561 & ~n_17364;
assign n_17368 = ~n_17363 &  n_17367;
assign n_17369 =  n_16932 & ~n_17368;
assign n_17370 = ~n_17366 &  n_17369;
assign n_17371 = ~n_17358 & ~n_17370;
assign n_17372 =  n_17346 &  n_17371;
assign n_17373 =  x_545 & ~n_17372;
assign n_17374 = ~x_545 &  n_17372;
assign n_17375 = ~n_17373 & ~n_17374;
assign n_17376 = ~x_1664 &  n_17328;
assign n_17377 =  x_1664 & ~n_17328;
assign n_17378 = ~n_17376 & ~n_17377;
assign n_17379 = ~n_17332 & ~n_17336;
assign n_17380 =  n_17378 & ~n_17379;
assign n_17381 = ~n_17378 &  n_17379;
assign n_17382 = ~n_17380 & ~n_17381;
assign n_17383 = ~x_288 & ~n_17382;
assign n_17384 =  x_288 & ~n_17381;
assign n_17385 = ~n_17380 &  n_17384;
assign n_17386 =  n_16927 & ~n_17385;
assign n_17387 = ~n_17383 &  n_17386;
assign n_17388 =  x_544 & ~n_16917;
assign n_17389 =  x_1024 & ~n_17342;
assign n_17390 = ~x_1024 &  n_17342;
assign n_17391 =  n_16925 & ~n_17390;
assign n_17392 = ~n_17389 &  n_17391;
assign n_17393 = ~n_17388 & ~n_17392;
assign n_17394 = ~n_17387 &  n_17393;
assign n_17395 = ~x_64 &  n_17347;
assign n_17396 =  x_64 & ~n_17347;
assign n_17397 = ~n_17395 & ~n_17396;
assign n_17398 = ~n_17351 & ~n_17355;
assign n_17399 =  n_17397 & ~n_17398;
assign n_17400 = ~n_17397 &  n_17398;
assign n_17401 = ~n_17399 & ~n_17400;
assign n_17402 = ~x_1952 & ~n_17401;
assign n_17403 =  x_1952 & ~n_17400;
assign n_17404 = ~n_17399 &  n_17403;
assign n_17405 =  n_16920 & ~n_17404;
assign n_17406 = ~n_17402 &  n_17405;
assign n_17407 = ~x_2624 &  n_17359;
assign n_17408 =  x_2624 & ~n_17359;
assign n_17409 = ~n_17407 & ~n_17408;
assign n_17410 = ~n_17363 & ~n_17367;
assign n_17411 =  n_17409 & ~n_17410;
assign n_17412 = ~n_17409 &  n_17410;
assign n_17413 = ~n_17411 & ~n_17412;
assign n_17414 = ~x_2560 & ~n_17413;
assign n_17415 =  x_2560 & ~n_17412;
assign n_17416 = ~n_17411 &  n_17415;
assign n_17417 =  n_16932 & ~n_17416;
assign n_17418 = ~n_17414 &  n_17417;
assign n_17419 = ~n_17406 & ~n_17418;
assign n_17420 =  n_17394 &  n_17419;
assign n_17421 =  x_544 & ~n_17420;
assign n_17422 = ~x_544 &  n_17420;
assign n_17423 = ~n_17421 & ~n_17422;
assign n_17424 = ~x_1663 &  n_17376;
assign n_17425 =  x_1663 & ~n_17376;
assign n_17426 = ~n_17424 & ~n_17425;
assign n_17427 = ~n_17380 & ~n_17384;
assign n_17428 =  n_17426 & ~n_17427;
assign n_17429 = ~n_17426 &  n_17427;
assign n_17430 = ~n_17428 & ~n_17429;
assign n_17431 = ~x_287 & ~n_17430;
assign n_17432 =  x_287 & ~n_17429;
assign n_17433 = ~n_17428 &  n_17432;
assign n_17434 =  n_16927 & ~n_17433;
assign n_17435 = ~n_17431 &  n_17434;
assign n_17436 =  x_543 & ~n_16917;
assign n_17437 =  x_1023 & ~n_17390;
assign n_17438 = ~x_1023 &  n_17390;
assign n_17439 =  n_16925 & ~n_17438;
assign n_17440 = ~n_17437 &  n_17439;
assign n_17441 = ~n_17436 & ~n_17440;
assign n_17442 = ~n_17435 &  n_17441;
assign n_17443 = ~x_63 &  n_17395;
assign n_17444 =  x_63 & ~n_17395;
assign n_17445 = ~n_17443 & ~n_17444;
assign n_17446 = ~n_17399 & ~n_17403;
assign n_17447 =  n_17445 & ~n_17446;
assign n_17448 = ~n_17445 &  n_17446;
assign n_17449 = ~n_17447 & ~n_17448;
assign n_17450 = ~x_1951 & ~n_17449;
assign n_17451 =  x_1951 & ~n_17448;
assign n_17452 = ~n_17447 &  n_17451;
assign n_17453 =  n_16920 & ~n_17452;
assign n_17454 = ~n_17450 &  n_17453;
assign n_17455 = ~x_2623 &  n_17407;
assign n_17456 =  x_2623 & ~n_17407;
assign n_17457 = ~n_17455 & ~n_17456;
assign n_17458 = ~n_17411 & ~n_17415;
assign n_17459 =  n_17457 & ~n_17458;
assign n_17460 = ~n_17457 &  n_17458;
assign n_17461 = ~n_17459 & ~n_17460;
assign n_17462 = ~x_2559 & ~n_17461;
assign n_17463 =  x_2559 & ~n_17460;
assign n_17464 = ~n_17459 &  n_17463;
assign n_17465 =  n_16932 & ~n_17464;
assign n_17466 = ~n_17462 &  n_17465;
assign n_17467 = ~n_17454 & ~n_17466;
assign n_17468 =  n_17442 &  n_17467;
assign n_17469 =  x_543 & ~n_17468;
assign n_17470 = ~x_543 &  n_17468;
assign n_17471 = ~n_17469 & ~n_17470;
assign n_17472 = ~x_1662 &  n_17424;
assign n_17473 =  x_1662 & ~n_17424;
assign n_17474 = ~n_17472 & ~n_17473;
assign n_17475 = ~n_17428 & ~n_17432;
assign n_17476 =  n_17474 & ~n_17475;
assign n_17477 = ~n_17474 &  n_17475;
assign n_17478 = ~n_17476 & ~n_17477;
assign n_17479 = ~x_286 & ~n_17478;
assign n_17480 =  x_286 & ~n_17477;
assign n_17481 = ~n_17476 &  n_17480;
assign n_17482 =  n_16927 & ~n_17481;
assign n_17483 = ~n_17479 &  n_17482;
assign n_17484 =  x_542 & ~n_16917;
assign n_17485 =  x_1022 & ~n_17438;
assign n_17486 = ~x_1022 &  n_17438;
assign n_17487 =  n_16925 & ~n_17486;
assign n_17488 = ~n_17485 &  n_17487;
assign n_17489 = ~n_17484 & ~n_17488;
assign n_17490 = ~n_17483 &  n_17489;
assign n_17491 = ~x_62 &  n_17443;
assign n_17492 =  x_62 & ~n_17443;
assign n_17493 = ~n_17491 & ~n_17492;
assign n_17494 = ~n_17447 & ~n_17451;
assign n_17495 =  n_17493 & ~n_17494;
assign n_17496 = ~n_17493 &  n_17494;
assign n_17497 = ~n_17495 & ~n_17496;
assign n_17498 = ~x_1950 & ~n_17497;
assign n_17499 =  x_1950 & ~n_17496;
assign n_17500 = ~n_17495 &  n_17499;
assign n_17501 =  n_16920 & ~n_17500;
assign n_17502 = ~n_17498 &  n_17501;
assign n_17503 = ~x_2622 &  n_17455;
assign n_17504 =  x_2622 & ~n_17455;
assign n_17505 = ~n_17503 & ~n_17504;
assign n_17506 = ~n_17459 & ~n_17463;
assign n_17507 =  n_17505 & ~n_17506;
assign n_17508 = ~n_17505 &  n_17506;
assign n_17509 = ~n_17507 & ~n_17508;
assign n_17510 = ~x_2558 & ~n_17509;
assign n_17511 =  x_2558 & ~n_17508;
assign n_17512 = ~n_17507 &  n_17511;
assign n_17513 =  n_16932 & ~n_17512;
assign n_17514 = ~n_17510 &  n_17513;
assign n_17515 = ~n_17502 & ~n_17514;
assign n_17516 =  n_17490 &  n_17515;
assign n_17517 =  x_542 & ~n_17516;
assign n_17518 = ~x_542 &  n_17516;
assign n_17519 = ~n_17517 & ~n_17518;
assign n_17520 = ~x_1661 &  n_17472;
assign n_17521 =  x_1661 & ~n_17472;
assign n_17522 = ~n_17520 & ~n_17521;
assign n_17523 = ~n_17476 & ~n_17480;
assign n_17524 =  n_17522 & ~n_17523;
assign n_17525 = ~n_17522 &  n_17523;
assign n_17526 = ~n_17524 & ~n_17525;
assign n_17527 = ~x_285 & ~n_17526;
assign n_17528 =  x_285 & ~n_17525;
assign n_17529 = ~n_17524 &  n_17528;
assign n_17530 =  n_16927 & ~n_17529;
assign n_17531 = ~n_17527 &  n_17530;
assign n_17532 =  x_541 & ~n_16917;
assign n_17533 =  x_1021 & ~n_17486;
assign n_17534 = ~x_1021 &  n_17486;
assign n_17535 =  n_16925 & ~n_17534;
assign n_17536 = ~n_17533 &  n_17535;
assign n_17537 = ~n_17532 & ~n_17536;
assign n_17538 = ~n_17531 &  n_17537;
assign n_17539 = ~x_61 &  n_17491;
assign n_17540 =  x_61 & ~n_17491;
assign n_17541 = ~n_17539 & ~n_17540;
assign n_17542 = ~n_17495 & ~n_17499;
assign n_17543 =  n_17541 & ~n_17542;
assign n_17544 = ~n_17541 &  n_17542;
assign n_17545 = ~n_17543 & ~n_17544;
assign n_17546 = ~x_1949 & ~n_17545;
assign n_17547 =  x_1949 & ~n_17544;
assign n_17548 = ~n_17543 &  n_17547;
assign n_17549 =  n_16920 & ~n_17548;
assign n_17550 = ~n_17546 &  n_17549;
assign n_17551 = ~x_2621 &  n_17503;
assign n_17552 =  x_2621 & ~n_17503;
assign n_17553 = ~n_17551 & ~n_17552;
assign n_17554 = ~n_17507 & ~n_17511;
assign n_17555 =  n_17553 & ~n_17554;
assign n_17556 = ~n_17553 &  n_17554;
assign n_17557 = ~n_17555 & ~n_17556;
assign n_17558 = ~x_2557 & ~n_17557;
assign n_17559 =  x_2557 & ~n_17556;
assign n_17560 = ~n_17555 &  n_17559;
assign n_17561 =  n_16932 & ~n_17560;
assign n_17562 = ~n_17558 &  n_17561;
assign n_17563 = ~n_17550 & ~n_17562;
assign n_17564 =  n_17538 &  n_17563;
assign n_17565 =  x_541 & ~n_17564;
assign n_17566 = ~x_541 &  n_17564;
assign n_17567 = ~n_17565 & ~n_17566;
assign n_17568 = ~x_1660 &  n_17520;
assign n_17569 =  x_1660 & ~n_17520;
assign n_17570 = ~n_17568 & ~n_17569;
assign n_17571 = ~n_17524 & ~n_17528;
assign n_17572 =  n_17570 & ~n_17571;
assign n_17573 = ~n_17570 &  n_17571;
assign n_17574 = ~n_17572 & ~n_17573;
assign n_17575 = ~x_284 & ~n_17574;
assign n_17576 =  x_284 & ~n_17573;
assign n_17577 = ~n_17572 &  n_17576;
assign n_17578 =  n_16927 & ~n_17577;
assign n_17579 = ~n_17575 &  n_17578;
assign n_17580 =  x_540 & ~n_16917;
assign n_17581 =  x_1020 & ~n_17534;
assign n_17582 = ~x_1020 &  n_17534;
assign n_17583 =  n_16925 & ~n_17582;
assign n_17584 = ~n_17581 &  n_17583;
assign n_17585 = ~n_17580 & ~n_17584;
assign n_17586 = ~n_17579 &  n_17585;
assign n_17587 = ~x_60 &  n_17539;
assign n_17588 =  x_60 & ~n_17539;
assign n_17589 = ~n_17587 & ~n_17588;
assign n_17590 = ~n_17543 & ~n_17547;
assign n_17591 =  n_17589 & ~n_17590;
assign n_17592 = ~n_17589 &  n_17590;
assign n_17593 = ~n_17591 & ~n_17592;
assign n_17594 = ~x_1948 & ~n_17593;
assign n_17595 =  x_1948 & ~n_17592;
assign n_17596 = ~n_17591 &  n_17595;
assign n_17597 =  n_16920 & ~n_17596;
assign n_17598 = ~n_17594 &  n_17597;
assign n_17599 = ~x_2620 &  n_17551;
assign n_17600 =  x_2620 & ~n_17551;
assign n_17601 = ~n_17599 & ~n_17600;
assign n_17602 = ~n_17555 & ~n_17559;
assign n_17603 =  n_17601 & ~n_17602;
assign n_17604 = ~n_17601 &  n_17602;
assign n_17605 = ~n_17603 & ~n_17604;
assign n_17606 = ~x_2556 & ~n_17605;
assign n_17607 =  x_2556 & ~n_17604;
assign n_17608 = ~n_17603 &  n_17607;
assign n_17609 =  n_16932 & ~n_17608;
assign n_17610 = ~n_17606 &  n_17609;
assign n_17611 = ~n_17598 & ~n_17610;
assign n_17612 =  n_17586 &  n_17611;
assign n_17613 =  x_540 & ~n_17612;
assign n_17614 = ~x_540 &  n_17612;
assign n_17615 = ~n_17613 & ~n_17614;
assign n_17616 = ~x_1659 &  n_17568;
assign n_17617 =  x_1659 & ~n_17568;
assign n_17618 = ~n_17616 & ~n_17617;
assign n_17619 = ~n_17572 & ~n_17576;
assign n_17620 =  n_17618 & ~n_17619;
assign n_17621 = ~n_17618 &  n_17619;
assign n_17622 = ~n_17620 & ~n_17621;
assign n_17623 = ~x_283 & ~n_17622;
assign n_17624 =  x_283 & ~n_17621;
assign n_17625 = ~n_17620 &  n_17624;
assign n_17626 =  n_16927 & ~n_17625;
assign n_17627 = ~n_17623 &  n_17626;
assign n_17628 =  x_539 & ~n_16917;
assign n_17629 =  x_1019 & ~n_17582;
assign n_17630 = ~x_1019 &  n_17582;
assign n_17631 =  n_16925 & ~n_17630;
assign n_17632 = ~n_17629 &  n_17631;
assign n_17633 = ~n_17628 & ~n_17632;
assign n_17634 = ~n_17627 &  n_17633;
assign n_17635 = ~x_59 &  n_17587;
assign n_17636 =  x_59 & ~n_17587;
assign n_17637 = ~n_17635 & ~n_17636;
assign n_17638 = ~n_17591 & ~n_17595;
assign n_17639 =  n_17637 & ~n_17638;
assign n_17640 = ~n_17637 &  n_17638;
assign n_17641 = ~n_17639 & ~n_17640;
assign n_17642 = ~x_1947 & ~n_17641;
assign n_17643 =  x_1947 & ~n_17640;
assign n_17644 = ~n_17639 &  n_17643;
assign n_17645 =  n_16920 & ~n_17644;
assign n_17646 = ~n_17642 &  n_17645;
assign n_17647 = ~x_2619 &  n_17599;
assign n_17648 =  x_2619 & ~n_17599;
assign n_17649 = ~n_17647 & ~n_17648;
assign n_17650 = ~n_17603 & ~n_17607;
assign n_17651 =  n_17649 & ~n_17650;
assign n_17652 = ~n_17649 &  n_17650;
assign n_17653 = ~n_17651 & ~n_17652;
assign n_17654 = ~x_2555 & ~n_17653;
assign n_17655 =  x_2555 & ~n_17652;
assign n_17656 = ~n_17651 &  n_17655;
assign n_17657 =  n_16932 & ~n_17656;
assign n_17658 = ~n_17654 &  n_17657;
assign n_17659 = ~n_17646 & ~n_17658;
assign n_17660 =  n_17634 &  n_17659;
assign n_17661 =  x_539 & ~n_17660;
assign n_17662 = ~x_539 &  n_17660;
assign n_17663 = ~n_17661 & ~n_17662;
assign n_17664 = ~x_1658 &  n_17616;
assign n_17665 =  x_1658 & ~n_17616;
assign n_17666 = ~n_17664 & ~n_17665;
assign n_17667 = ~n_17620 & ~n_17624;
assign n_17668 =  n_17666 & ~n_17667;
assign n_17669 = ~n_17666 &  n_17667;
assign n_17670 = ~n_17668 & ~n_17669;
assign n_17671 = ~x_282 & ~n_17670;
assign n_17672 =  x_282 & ~n_17669;
assign n_17673 = ~n_17668 &  n_17672;
assign n_17674 =  n_16927 & ~n_17673;
assign n_17675 = ~n_17671 &  n_17674;
assign n_17676 =  x_538 & ~n_16917;
assign n_17677 =  x_1018 & ~n_17630;
assign n_17678 = ~x_1018 &  n_17630;
assign n_17679 =  n_16925 & ~n_17678;
assign n_17680 = ~n_17677 &  n_17679;
assign n_17681 = ~n_17676 & ~n_17680;
assign n_17682 = ~n_17675 &  n_17681;
assign n_17683 = ~x_58 &  n_17635;
assign n_17684 =  x_58 & ~n_17635;
assign n_17685 = ~n_17683 & ~n_17684;
assign n_17686 = ~n_17639 & ~n_17643;
assign n_17687 =  n_17685 & ~n_17686;
assign n_17688 = ~n_17685 &  n_17686;
assign n_17689 = ~n_17687 & ~n_17688;
assign n_17690 = ~x_1946 & ~n_17689;
assign n_17691 =  x_1946 & ~n_17688;
assign n_17692 = ~n_17687 &  n_17691;
assign n_17693 =  n_16920 & ~n_17692;
assign n_17694 = ~n_17690 &  n_17693;
assign n_17695 = ~x_2618 &  n_17647;
assign n_17696 =  x_2618 & ~n_17647;
assign n_17697 = ~n_17695 & ~n_17696;
assign n_17698 = ~n_17651 & ~n_17655;
assign n_17699 =  n_17697 & ~n_17698;
assign n_17700 = ~n_17697 &  n_17698;
assign n_17701 = ~n_17699 & ~n_17700;
assign n_17702 = ~x_2554 & ~n_17701;
assign n_17703 =  x_2554 & ~n_17700;
assign n_17704 = ~n_17699 &  n_17703;
assign n_17705 =  n_16932 & ~n_17704;
assign n_17706 = ~n_17702 &  n_17705;
assign n_17707 = ~n_17694 & ~n_17706;
assign n_17708 =  n_17682 &  n_17707;
assign n_17709 =  x_538 & ~n_17708;
assign n_17710 = ~x_538 &  n_17708;
assign n_17711 = ~n_17709 & ~n_17710;
assign n_17712 = ~x_1657 &  n_17664;
assign n_17713 =  x_1657 & ~n_17664;
assign n_17714 = ~n_17712 & ~n_17713;
assign n_17715 = ~n_17668 & ~n_17672;
assign n_17716 =  n_17714 & ~n_17715;
assign n_17717 = ~n_17714 &  n_17715;
assign n_17718 = ~n_17716 & ~n_17717;
assign n_17719 = ~x_281 & ~n_17718;
assign n_17720 =  x_281 & ~n_17717;
assign n_17721 = ~n_17716 &  n_17720;
assign n_17722 =  n_16927 & ~n_17721;
assign n_17723 = ~n_17719 &  n_17722;
assign n_17724 =  x_537 & ~n_16917;
assign n_17725 =  x_1017 & ~n_17678;
assign n_17726 = ~x_1017 &  n_17678;
assign n_17727 =  n_16925 & ~n_17726;
assign n_17728 = ~n_17725 &  n_17727;
assign n_17729 = ~n_17724 & ~n_17728;
assign n_17730 = ~n_17723 &  n_17729;
assign n_17731 = ~x_57 &  n_17683;
assign n_17732 =  x_57 & ~n_17683;
assign n_17733 = ~n_17731 & ~n_17732;
assign n_17734 = ~n_17687 & ~n_17691;
assign n_17735 =  n_17733 & ~n_17734;
assign n_17736 = ~n_17733 &  n_17734;
assign n_17737 = ~n_17735 & ~n_17736;
assign n_17738 = ~x_1945 & ~n_17737;
assign n_17739 =  x_1945 & ~n_17736;
assign n_17740 = ~n_17735 &  n_17739;
assign n_17741 =  n_16920 & ~n_17740;
assign n_17742 = ~n_17738 &  n_17741;
assign n_17743 = ~x_2617 &  n_17695;
assign n_17744 =  x_2617 & ~n_17695;
assign n_17745 = ~n_17743 & ~n_17744;
assign n_17746 = ~n_17699 & ~n_17703;
assign n_17747 =  n_17745 & ~n_17746;
assign n_17748 = ~n_17745 &  n_17746;
assign n_17749 = ~n_17747 & ~n_17748;
assign n_17750 = ~x_2553 & ~n_17749;
assign n_17751 =  x_2553 & ~n_17748;
assign n_17752 = ~n_17747 &  n_17751;
assign n_17753 =  n_16932 & ~n_17752;
assign n_17754 = ~n_17750 &  n_17753;
assign n_17755 = ~n_17742 & ~n_17754;
assign n_17756 =  n_17730 &  n_17755;
assign n_17757 =  x_537 & ~n_17756;
assign n_17758 = ~x_537 &  n_17756;
assign n_17759 = ~n_17757 & ~n_17758;
assign n_17760 = ~x_1656 &  n_17712;
assign n_17761 =  x_1656 & ~n_17712;
assign n_17762 = ~n_17760 & ~n_17761;
assign n_17763 = ~n_17716 & ~n_17720;
assign n_17764 =  n_17762 & ~n_17763;
assign n_17765 = ~n_17762 &  n_17763;
assign n_17766 = ~n_17764 & ~n_17765;
assign n_17767 = ~x_280 & ~n_17766;
assign n_17768 =  x_280 & ~n_17765;
assign n_17769 = ~n_17764 &  n_17768;
assign n_17770 =  n_16927 & ~n_17769;
assign n_17771 = ~n_17767 &  n_17770;
assign n_17772 =  x_536 & ~n_16917;
assign n_17773 =  x_1016 & ~n_17726;
assign n_17774 = ~x_1016 &  n_17726;
assign n_17775 =  n_16925 & ~n_17774;
assign n_17776 = ~n_17773 &  n_17775;
assign n_17777 = ~n_17772 & ~n_17776;
assign n_17778 = ~n_17771 &  n_17777;
assign n_17779 = ~x_56 &  n_17731;
assign n_17780 =  x_56 & ~n_17731;
assign n_17781 = ~n_17779 & ~n_17780;
assign n_17782 = ~n_17735 & ~n_17739;
assign n_17783 =  n_17781 & ~n_17782;
assign n_17784 = ~n_17781 &  n_17782;
assign n_17785 = ~n_17783 & ~n_17784;
assign n_17786 = ~x_1944 & ~n_17785;
assign n_17787 =  x_1944 & ~n_17784;
assign n_17788 = ~n_17783 &  n_17787;
assign n_17789 =  n_16920 & ~n_17788;
assign n_17790 = ~n_17786 &  n_17789;
assign n_17791 = ~x_2616 &  n_17743;
assign n_17792 =  x_2616 & ~n_17743;
assign n_17793 = ~n_17791 & ~n_17792;
assign n_17794 = ~n_17747 & ~n_17751;
assign n_17795 =  n_17793 & ~n_17794;
assign n_17796 = ~n_17793 &  n_17794;
assign n_17797 = ~n_17795 & ~n_17796;
assign n_17798 = ~x_2552 & ~n_17797;
assign n_17799 =  x_2552 & ~n_17796;
assign n_17800 = ~n_17795 &  n_17799;
assign n_17801 =  n_16932 & ~n_17800;
assign n_17802 = ~n_17798 &  n_17801;
assign n_17803 = ~n_17790 & ~n_17802;
assign n_17804 =  n_17778 &  n_17803;
assign n_17805 =  x_536 & ~n_17804;
assign n_17806 = ~x_536 &  n_17804;
assign n_17807 = ~n_17805 & ~n_17806;
assign n_17808 = ~x_1655 &  n_17760;
assign n_17809 =  x_1655 & ~n_17760;
assign n_17810 = ~n_17808 & ~n_17809;
assign n_17811 = ~n_17764 & ~n_17768;
assign n_17812 =  n_17810 & ~n_17811;
assign n_17813 = ~n_17810 &  n_17811;
assign n_17814 = ~n_17812 & ~n_17813;
assign n_17815 = ~x_279 & ~n_17814;
assign n_17816 =  x_279 & ~n_17813;
assign n_17817 = ~n_17812 &  n_17816;
assign n_17818 =  n_16927 & ~n_17817;
assign n_17819 = ~n_17815 &  n_17818;
assign n_17820 =  x_535 & ~n_16917;
assign n_17821 =  x_1015 & ~n_17774;
assign n_17822 = ~x_1015 &  n_17774;
assign n_17823 =  n_16925 & ~n_17822;
assign n_17824 = ~n_17821 &  n_17823;
assign n_17825 = ~n_17820 & ~n_17824;
assign n_17826 = ~n_17819 &  n_17825;
assign n_17827 = ~x_55 &  n_17779;
assign n_17828 =  x_55 & ~n_17779;
assign n_17829 = ~n_17827 & ~n_17828;
assign n_17830 = ~n_17783 & ~n_17787;
assign n_17831 =  n_17829 & ~n_17830;
assign n_17832 = ~n_17829 &  n_17830;
assign n_17833 = ~n_17831 & ~n_17832;
assign n_17834 = ~x_1943 & ~n_17833;
assign n_17835 =  x_1943 & ~n_17832;
assign n_17836 = ~n_17831 &  n_17835;
assign n_17837 =  n_16920 & ~n_17836;
assign n_17838 = ~n_17834 &  n_17837;
assign n_17839 = ~x_2615 &  n_17791;
assign n_17840 =  x_2615 & ~n_17791;
assign n_17841 = ~n_17839 & ~n_17840;
assign n_17842 = ~n_17795 & ~n_17799;
assign n_17843 =  n_17841 & ~n_17842;
assign n_17844 = ~n_17841 &  n_17842;
assign n_17845 = ~n_17843 & ~n_17844;
assign n_17846 = ~x_2551 & ~n_17845;
assign n_17847 =  x_2551 & ~n_17844;
assign n_17848 = ~n_17843 &  n_17847;
assign n_17849 =  n_16932 & ~n_17848;
assign n_17850 = ~n_17846 &  n_17849;
assign n_17851 = ~n_17838 & ~n_17850;
assign n_17852 =  n_17826 &  n_17851;
assign n_17853 =  x_535 & ~n_17852;
assign n_17854 = ~x_535 &  n_17852;
assign n_17855 = ~n_17853 & ~n_17854;
assign n_17856 = ~x_1654 &  n_17808;
assign n_17857 =  x_1654 & ~n_17808;
assign n_17858 = ~n_17856 & ~n_17857;
assign n_17859 = ~n_17812 & ~n_17816;
assign n_17860 =  n_17858 & ~n_17859;
assign n_17861 = ~n_17858 &  n_17859;
assign n_17862 = ~n_17860 & ~n_17861;
assign n_17863 = ~x_278 & ~n_17862;
assign n_17864 =  x_278 & ~n_17861;
assign n_17865 = ~n_17860 &  n_17864;
assign n_17866 =  n_16927 & ~n_17865;
assign n_17867 = ~n_17863 &  n_17866;
assign n_17868 =  x_534 & ~n_16917;
assign n_17869 =  x_1014 & ~n_17822;
assign n_17870 = ~x_1014 &  n_17822;
assign n_17871 =  n_16925 & ~n_17870;
assign n_17872 = ~n_17869 &  n_17871;
assign n_17873 = ~n_17868 & ~n_17872;
assign n_17874 = ~n_17867 &  n_17873;
assign n_17875 = ~x_54 &  n_17827;
assign n_17876 =  x_54 & ~n_17827;
assign n_17877 = ~n_17875 & ~n_17876;
assign n_17878 = ~n_17831 & ~n_17835;
assign n_17879 =  n_17877 & ~n_17878;
assign n_17880 = ~n_17877 &  n_17878;
assign n_17881 = ~n_17879 & ~n_17880;
assign n_17882 = ~x_1942 & ~n_17881;
assign n_17883 =  x_1942 & ~n_17880;
assign n_17884 = ~n_17879 &  n_17883;
assign n_17885 =  n_16920 & ~n_17884;
assign n_17886 = ~n_17882 &  n_17885;
assign n_17887 = ~x_2614 &  n_17839;
assign n_17888 =  x_2614 & ~n_17839;
assign n_17889 = ~n_17887 & ~n_17888;
assign n_17890 = ~n_17843 & ~n_17847;
assign n_17891 =  n_17889 & ~n_17890;
assign n_17892 = ~n_17889 &  n_17890;
assign n_17893 = ~n_17891 & ~n_17892;
assign n_17894 = ~x_2550 & ~n_17893;
assign n_17895 =  x_2550 & ~n_17892;
assign n_17896 = ~n_17891 &  n_17895;
assign n_17897 =  n_16932 & ~n_17896;
assign n_17898 = ~n_17894 &  n_17897;
assign n_17899 = ~n_17886 & ~n_17898;
assign n_17900 =  n_17874 &  n_17899;
assign n_17901 =  x_534 & ~n_17900;
assign n_17902 = ~x_534 &  n_17900;
assign n_17903 = ~n_17901 & ~n_17902;
assign n_17904 = ~x_1653 &  n_17856;
assign n_17905 =  x_1653 & ~n_17856;
assign n_17906 = ~n_17904 & ~n_17905;
assign n_17907 = ~n_17860 & ~n_17864;
assign n_17908 =  n_17906 & ~n_17907;
assign n_17909 = ~n_17906 &  n_17907;
assign n_17910 = ~n_17908 & ~n_17909;
assign n_17911 = ~x_277 & ~n_17910;
assign n_17912 =  x_277 & ~n_17909;
assign n_17913 = ~n_17908 &  n_17912;
assign n_17914 =  n_16927 & ~n_17913;
assign n_17915 = ~n_17911 &  n_17914;
assign n_17916 =  x_533 & ~n_16917;
assign n_17917 =  x_1013 & ~n_17870;
assign n_17918 = ~x_1013 &  n_17870;
assign n_17919 =  n_16925 & ~n_17918;
assign n_17920 = ~n_17917 &  n_17919;
assign n_17921 = ~n_17916 & ~n_17920;
assign n_17922 = ~n_17915 &  n_17921;
assign n_17923 = ~x_53 &  n_17875;
assign n_17924 =  x_53 & ~n_17875;
assign n_17925 = ~n_17923 & ~n_17924;
assign n_17926 = ~n_17879 & ~n_17883;
assign n_17927 =  n_17925 & ~n_17926;
assign n_17928 = ~n_17925 &  n_17926;
assign n_17929 = ~n_17927 & ~n_17928;
assign n_17930 = ~x_1941 & ~n_17929;
assign n_17931 =  x_1941 & ~n_17928;
assign n_17932 = ~n_17927 &  n_17931;
assign n_17933 =  n_16920 & ~n_17932;
assign n_17934 = ~n_17930 &  n_17933;
assign n_17935 = ~x_2613 &  n_17887;
assign n_17936 =  x_2613 & ~n_17887;
assign n_17937 = ~n_17935 & ~n_17936;
assign n_17938 = ~n_17891 & ~n_17895;
assign n_17939 =  n_17937 & ~n_17938;
assign n_17940 = ~n_17937 &  n_17938;
assign n_17941 = ~n_17939 & ~n_17940;
assign n_17942 = ~x_2549 & ~n_17941;
assign n_17943 =  x_2549 & ~n_17940;
assign n_17944 = ~n_17939 &  n_17943;
assign n_17945 =  n_16932 & ~n_17944;
assign n_17946 = ~n_17942 &  n_17945;
assign n_17947 = ~n_17934 & ~n_17946;
assign n_17948 =  n_17922 &  n_17947;
assign n_17949 =  x_533 & ~n_17948;
assign n_17950 = ~x_533 &  n_17948;
assign n_17951 = ~n_17949 & ~n_17950;
assign n_17952 = ~x_1652 &  n_17904;
assign n_17953 =  x_1652 & ~n_17904;
assign n_17954 = ~n_17952 & ~n_17953;
assign n_17955 = ~n_17908 & ~n_17912;
assign n_17956 =  n_17954 & ~n_17955;
assign n_17957 = ~n_17954 &  n_17955;
assign n_17958 = ~n_17956 & ~n_17957;
assign n_17959 = ~x_276 & ~n_17958;
assign n_17960 =  x_276 & ~n_17957;
assign n_17961 = ~n_17956 &  n_17960;
assign n_17962 =  n_16927 & ~n_17961;
assign n_17963 = ~n_17959 &  n_17962;
assign n_17964 =  x_532 & ~n_16917;
assign n_17965 =  x_1012 & ~n_17918;
assign n_17966 = ~x_1012 &  n_17918;
assign n_17967 =  n_16925 & ~n_17966;
assign n_17968 = ~n_17965 &  n_17967;
assign n_17969 = ~n_17964 & ~n_17968;
assign n_17970 = ~n_17963 &  n_17969;
assign n_17971 = ~x_52 &  n_17923;
assign n_17972 =  x_52 & ~n_17923;
assign n_17973 = ~n_17971 & ~n_17972;
assign n_17974 = ~n_17927 & ~n_17931;
assign n_17975 =  n_17973 & ~n_17974;
assign n_17976 = ~n_17973 &  n_17974;
assign n_17977 = ~n_17975 & ~n_17976;
assign n_17978 = ~x_1940 & ~n_17977;
assign n_17979 =  x_1940 & ~n_17976;
assign n_17980 = ~n_17975 &  n_17979;
assign n_17981 =  n_16920 & ~n_17980;
assign n_17982 = ~n_17978 &  n_17981;
assign n_17983 = ~x_2612 &  n_17935;
assign n_17984 =  x_2612 & ~n_17935;
assign n_17985 = ~n_17983 & ~n_17984;
assign n_17986 = ~n_17939 & ~n_17943;
assign n_17987 =  n_17985 & ~n_17986;
assign n_17988 = ~n_17985 &  n_17986;
assign n_17989 = ~n_17987 & ~n_17988;
assign n_17990 = ~x_2548 & ~n_17989;
assign n_17991 =  x_2548 & ~n_17988;
assign n_17992 = ~n_17987 &  n_17991;
assign n_17993 =  n_16932 & ~n_17992;
assign n_17994 = ~n_17990 &  n_17993;
assign n_17995 = ~n_17982 & ~n_17994;
assign n_17996 =  n_17970 &  n_17995;
assign n_17997 =  x_532 & ~n_17996;
assign n_17998 = ~x_532 &  n_17996;
assign n_17999 = ~n_17997 & ~n_17998;
assign n_18000 = ~x_1651 &  n_17952;
assign n_18001 =  x_1651 & ~n_17952;
assign n_18002 = ~n_18000 & ~n_18001;
assign n_18003 = ~n_17956 & ~n_17960;
assign n_18004 =  n_18002 & ~n_18003;
assign n_18005 = ~n_18002 &  n_18003;
assign n_18006 = ~n_18004 & ~n_18005;
assign n_18007 = ~x_275 & ~n_18006;
assign n_18008 =  x_275 & ~n_18005;
assign n_18009 = ~n_18004 &  n_18008;
assign n_18010 =  n_16927 & ~n_18009;
assign n_18011 = ~n_18007 &  n_18010;
assign n_18012 =  x_531 & ~n_16917;
assign n_18013 =  x_1011 & ~n_17966;
assign n_18014 = ~x_1011 &  n_17966;
assign n_18015 =  n_16925 & ~n_18014;
assign n_18016 = ~n_18013 &  n_18015;
assign n_18017 = ~n_18012 & ~n_18016;
assign n_18018 = ~n_18011 &  n_18017;
assign n_18019 = ~x_51 &  n_17971;
assign n_18020 =  x_51 & ~n_17971;
assign n_18021 = ~n_18019 & ~n_18020;
assign n_18022 = ~n_17975 & ~n_17979;
assign n_18023 =  n_18021 & ~n_18022;
assign n_18024 = ~n_18021 &  n_18022;
assign n_18025 = ~n_18023 & ~n_18024;
assign n_18026 = ~x_1939 & ~n_18025;
assign n_18027 =  x_1939 & ~n_18024;
assign n_18028 = ~n_18023 &  n_18027;
assign n_18029 =  n_16920 & ~n_18028;
assign n_18030 = ~n_18026 &  n_18029;
assign n_18031 = ~x_2611 &  n_17983;
assign n_18032 =  x_2611 & ~n_17983;
assign n_18033 = ~n_18031 & ~n_18032;
assign n_18034 = ~n_17987 & ~n_17991;
assign n_18035 =  n_18033 & ~n_18034;
assign n_18036 = ~n_18033 &  n_18034;
assign n_18037 = ~n_18035 & ~n_18036;
assign n_18038 = ~x_2547 & ~n_18037;
assign n_18039 =  x_2547 & ~n_18036;
assign n_18040 = ~n_18035 &  n_18039;
assign n_18041 =  n_16932 & ~n_18040;
assign n_18042 = ~n_18038 &  n_18041;
assign n_18043 = ~n_18030 & ~n_18042;
assign n_18044 =  n_18018 &  n_18043;
assign n_18045 =  x_531 & ~n_18044;
assign n_18046 = ~x_531 &  n_18044;
assign n_18047 = ~n_18045 & ~n_18046;
assign n_18048 = ~x_1650 &  n_18000;
assign n_18049 =  x_1650 & ~n_18000;
assign n_18050 = ~n_18048 & ~n_18049;
assign n_18051 = ~n_18004 & ~n_18008;
assign n_18052 =  n_18050 & ~n_18051;
assign n_18053 = ~n_18050 &  n_18051;
assign n_18054 = ~n_18052 & ~n_18053;
assign n_18055 = ~x_274 & ~n_18054;
assign n_18056 =  x_274 & ~n_18053;
assign n_18057 = ~n_18052 &  n_18056;
assign n_18058 =  n_16927 & ~n_18057;
assign n_18059 = ~n_18055 &  n_18058;
assign n_18060 =  x_530 & ~n_16917;
assign n_18061 =  x_1010 & ~n_18014;
assign n_18062 = ~x_1010 &  n_18014;
assign n_18063 =  n_16925 & ~n_18062;
assign n_18064 = ~n_18061 &  n_18063;
assign n_18065 = ~n_18060 & ~n_18064;
assign n_18066 = ~n_18059 &  n_18065;
assign n_18067 = ~x_50 &  n_18019;
assign n_18068 =  x_50 & ~n_18019;
assign n_18069 = ~n_18067 & ~n_18068;
assign n_18070 = ~n_18023 & ~n_18027;
assign n_18071 =  n_18069 & ~n_18070;
assign n_18072 = ~n_18069 &  n_18070;
assign n_18073 = ~n_18071 & ~n_18072;
assign n_18074 = ~x_1938 & ~n_18073;
assign n_18075 =  x_1938 & ~n_18072;
assign n_18076 = ~n_18071 &  n_18075;
assign n_18077 =  n_16920 & ~n_18076;
assign n_18078 = ~n_18074 &  n_18077;
assign n_18079 = ~x_2610 &  n_18031;
assign n_18080 =  x_2610 & ~n_18031;
assign n_18081 = ~n_18079 & ~n_18080;
assign n_18082 = ~n_18035 & ~n_18039;
assign n_18083 =  n_18081 & ~n_18082;
assign n_18084 = ~n_18081 &  n_18082;
assign n_18085 = ~n_18083 & ~n_18084;
assign n_18086 = ~x_2546 & ~n_18085;
assign n_18087 =  x_2546 & ~n_18084;
assign n_18088 = ~n_18083 &  n_18087;
assign n_18089 =  n_16932 & ~n_18088;
assign n_18090 = ~n_18086 &  n_18089;
assign n_18091 = ~n_18078 & ~n_18090;
assign n_18092 =  n_18066 &  n_18091;
assign n_18093 =  x_530 & ~n_18092;
assign n_18094 = ~x_530 &  n_18092;
assign n_18095 = ~n_18093 & ~n_18094;
assign n_18096 = ~x_1649 &  n_18048;
assign n_18097 =  x_1649 & ~n_18048;
assign n_18098 = ~n_18096 & ~n_18097;
assign n_18099 = ~n_18052 & ~n_18056;
assign n_18100 =  n_18098 & ~n_18099;
assign n_18101 = ~n_18098 &  n_18099;
assign n_18102 = ~n_18100 & ~n_18101;
assign n_18103 = ~x_273 & ~n_18102;
assign n_18104 =  x_273 & ~n_18101;
assign n_18105 = ~n_18100 &  n_18104;
assign n_18106 =  n_16927 & ~n_18105;
assign n_18107 = ~n_18103 &  n_18106;
assign n_18108 =  x_529 & ~n_16917;
assign n_18109 =  x_1009 & ~n_18062;
assign n_18110 = ~x_1009 &  n_18062;
assign n_18111 =  n_16925 & ~n_18110;
assign n_18112 = ~n_18109 &  n_18111;
assign n_18113 = ~n_18108 & ~n_18112;
assign n_18114 = ~n_18107 &  n_18113;
assign n_18115 = ~x_49 &  n_18067;
assign n_18116 =  x_49 & ~n_18067;
assign n_18117 = ~n_18115 & ~n_18116;
assign n_18118 = ~n_18071 & ~n_18075;
assign n_18119 =  n_18117 & ~n_18118;
assign n_18120 = ~n_18117 &  n_18118;
assign n_18121 = ~n_18119 & ~n_18120;
assign n_18122 = ~x_1937 & ~n_18121;
assign n_18123 =  x_1937 & ~n_18120;
assign n_18124 = ~n_18119 &  n_18123;
assign n_18125 =  n_16920 & ~n_18124;
assign n_18126 = ~n_18122 &  n_18125;
assign n_18127 = ~x_2609 &  n_18079;
assign n_18128 =  x_2609 & ~n_18079;
assign n_18129 = ~n_18127 & ~n_18128;
assign n_18130 = ~n_18083 & ~n_18087;
assign n_18131 =  n_18129 & ~n_18130;
assign n_18132 = ~n_18129 &  n_18130;
assign n_18133 = ~n_18131 & ~n_18132;
assign n_18134 = ~x_2545 & ~n_18133;
assign n_18135 =  x_2545 & ~n_18132;
assign n_18136 = ~n_18131 &  n_18135;
assign n_18137 =  n_16932 & ~n_18136;
assign n_18138 = ~n_18134 &  n_18137;
assign n_18139 = ~n_18126 & ~n_18138;
assign n_18140 =  n_18114 &  n_18139;
assign n_18141 =  x_529 & ~n_18140;
assign n_18142 = ~x_529 &  n_18140;
assign n_18143 = ~n_18141 & ~n_18142;
assign n_18144 = ~x_1648 &  n_18096;
assign n_18145 =  x_1648 & ~n_18096;
assign n_18146 = ~n_18144 & ~n_18145;
assign n_18147 = ~n_18100 & ~n_18104;
assign n_18148 =  n_18146 & ~n_18147;
assign n_18149 = ~n_18146 &  n_18147;
assign n_18150 = ~n_18148 & ~n_18149;
assign n_18151 = ~x_272 & ~n_18150;
assign n_18152 =  x_272 & ~n_18149;
assign n_18153 = ~n_18148 &  n_18152;
assign n_18154 =  n_16927 & ~n_18153;
assign n_18155 = ~n_18151 &  n_18154;
assign n_18156 =  x_528 & ~n_16917;
assign n_18157 =  x_1008 & ~n_18110;
assign n_18158 = ~x_1008 &  n_18110;
assign n_18159 =  n_16925 & ~n_18158;
assign n_18160 = ~n_18157 &  n_18159;
assign n_18161 = ~n_18156 & ~n_18160;
assign n_18162 = ~n_18155 &  n_18161;
assign n_18163 = ~x_48 &  n_18115;
assign n_18164 =  x_48 & ~n_18115;
assign n_18165 = ~n_18163 & ~n_18164;
assign n_18166 = ~n_18119 & ~n_18123;
assign n_18167 =  n_18165 & ~n_18166;
assign n_18168 = ~n_18165 &  n_18166;
assign n_18169 = ~n_18167 & ~n_18168;
assign n_18170 = ~x_1936 & ~n_18169;
assign n_18171 =  x_1936 & ~n_18168;
assign n_18172 = ~n_18167 &  n_18171;
assign n_18173 =  n_16920 & ~n_18172;
assign n_18174 = ~n_18170 &  n_18173;
assign n_18175 = ~x_2608 &  n_18127;
assign n_18176 =  x_2608 & ~n_18127;
assign n_18177 = ~n_18175 & ~n_18176;
assign n_18178 = ~n_18131 & ~n_18135;
assign n_18179 =  n_18177 & ~n_18178;
assign n_18180 = ~n_18177 &  n_18178;
assign n_18181 = ~n_18179 & ~n_18180;
assign n_18182 = ~x_2544 & ~n_18181;
assign n_18183 =  x_2544 & ~n_18180;
assign n_18184 = ~n_18179 &  n_18183;
assign n_18185 =  n_16932 & ~n_18184;
assign n_18186 = ~n_18182 &  n_18185;
assign n_18187 = ~n_18174 & ~n_18186;
assign n_18188 =  n_18162 &  n_18187;
assign n_18189 =  x_528 & ~n_18188;
assign n_18190 = ~x_528 &  n_18188;
assign n_18191 = ~n_18189 & ~n_18190;
assign n_18192 = ~x_1647 &  n_18144;
assign n_18193 =  x_1647 & ~n_18144;
assign n_18194 = ~n_18192 & ~n_18193;
assign n_18195 = ~n_18148 & ~n_18152;
assign n_18196 =  n_18194 & ~n_18195;
assign n_18197 = ~n_18194 &  n_18195;
assign n_18198 = ~n_18196 & ~n_18197;
assign n_18199 = ~x_271 & ~n_18198;
assign n_18200 =  x_271 & ~n_18197;
assign n_18201 = ~n_18196 &  n_18200;
assign n_18202 =  n_16927 & ~n_18201;
assign n_18203 = ~n_18199 &  n_18202;
assign n_18204 =  x_527 & ~n_16917;
assign n_18205 =  x_1007 & ~n_18158;
assign n_18206 = ~x_1007 &  n_18158;
assign n_18207 =  n_16925 & ~n_18206;
assign n_18208 = ~n_18205 &  n_18207;
assign n_18209 = ~n_18204 & ~n_18208;
assign n_18210 = ~n_18203 &  n_18209;
assign n_18211 = ~x_47 &  n_18163;
assign n_18212 =  x_47 & ~n_18163;
assign n_18213 = ~n_18211 & ~n_18212;
assign n_18214 = ~n_18167 & ~n_18171;
assign n_18215 =  n_18213 & ~n_18214;
assign n_18216 = ~n_18213 &  n_18214;
assign n_18217 = ~n_18215 & ~n_18216;
assign n_18218 = ~x_1935 & ~n_18217;
assign n_18219 =  x_1935 & ~n_18216;
assign n_18220 = ~n_18215 &  n_18219;
assign n_18221 =  n_16920 & ~n_18220;
assign n_18222 = ~n_18218 &  n_18221;
assign n_18223 = ~x_2607 &  n_18175;
assign n_18224 =  x_2607 & ~n_18175;
assign n_18225 = ~n_18223 & ~n_18224;
assign n_18226 = ~n_18179 & ~n_18183;
assign n_18227 =  n_18225 & ~n_18226;
assign n_18228 = ~n_18225 &  n_18226;
assign n_18229 = ~n_18227 & ~n_18228;
assign n_18230 = ~x_2543 & ~n_18229;
assign n_18231 =  x_2543 & ~n_18228;
assign n_18232 = ~n_18227 &  n_18231;
assign n_18233 =  n_16932 & ~n_18232;
assign n_18234 = ~n_18230 &  n_18233;
assign n_18235 = ~n_18222 & ~n_18234;
assign n_18236 =  n_18210 &  n_18235;
assign n_18237 =  x_527 & ~n_18236;
assign n_18238 = ~x_527 &  n_18236;
assign n_18239 = ~n_18237 & ~n_18238;
assign n_18240 = ~x_1646 &  n_18192;
assign n_18241 =  x_1646 & ~n_18192;
assign n_18242 = ~n_18240 & ~n_18241;
assign n_18243 = ~n_18196 & ~n_18200;
assign n_18244 =  n_18242 & ~n_18243;
assign n_18245 = ~n_18242 &  n_18243;
assign n_18246 = ~n_18244 & ~n_18245;
assign n_18247 = ~x_270 & ~n_18246;
assign n_18248 =  x_270 & ~n_18245;
assign n_18249 = ~n_18244 &  n_18248;
assign n_18250 =  n_16927 & ~n_18249;
assign n_18251 = ~n_18247 &  n_18250;
assign n_18252 =  x_526 & ~n_16917;
assign n_18253 =  x_1006 & ~n_18206;
assign n_18254 = ~x_1006 &  n_18206;
assign n_18255 =  n_16925 & ~n_18254;
assign n_18256 = ~n_18253 &  n_18255;
assign n_18257 = ~n_18252 & ~n_18256;
assign n_18258 = ~n_18251 &  n_18257;
assign n_18259 = ~x_46 &  n_18211;
assign n_18260 =  x_46 & ~n_18211;
assign n_18261 = ~n_18259 & ~n_18260;
assign n_18262 = ~n_18215 & ~n_18219;
assign n_18263 =  n_18261 & ~n_18262;
assign n_18264 = ~n_18261 &  n_18262;
assign n_18265 = ~n_18263 & ~n_18264;
assign n_18266 = ~x_1934 & ~n_18265;
assign n_18267 =  x_1934 & ~n_18264;
assign n_18268 = ~n_18263 &  n_18267;
assign n_18269 =  n_16920 & ~n_18268;
assign n_18270 = ~n_18266 &  n_18269;
assign n_18271 = ~x_2606 &  n_18223;
assign n_18272 =  x_2606 & ~n_18223;
assign n_18273 = ~n_18271 & ~n_18272;
assign n_18274 = ~n_18227 & ~n_18231;
assign n_18275 =  n_18273 & ~n_18274;
assign n_18276 = ~n_18273 &  n_18274;
assign n_18277 = ~n_18275 & ~n_18276;
assign n_18278 = ~x_2542 & ~n_18277;
assign n_18279 =  x_2542 & ~n_18276;
assign n_18280 = ~n_18275 &  n_18279;
assign n_18281 =  n_16932 & ~n_18280;
assign n_18282 = ~n_18278 &  n_18281;
assign n_18283 = ~n_18270 & ~n_18282;
assign n_18284 =  n_18258 &  n_18283;
assign n_18285 =  x_526 & ~n_18284;
assign n_18286 = ~x_526 &  n_18284;
assign n_18287 = ~n_18285 & ~n_18286;
assign n_18288 = ~x_1645 &  n_18240;
assign n_18289 =  x_1645 & ~n_18240;
assign n_18290 = ~n_18288 & ~n_18289;
assign n_18291 = ~n_18244 & ~n_18248;
assign n_18292 =  n_18290 & ~n_18291;
assign n_18293 = ~n_18290 &  n_18291;
assign n_18294 = ~n_18292 & ~n_18293;
assign n_18295 = ~x_269 & ~n_18294;
assign n_18296 =  x_269 & ~n_18293;
assign n_18297 = ~n_18292 &  n_18296;
assign n_18298 =  n_16927 & ~n_18297;
assign n_18299 = ~n_18295 &  n_18298;
assign n_18300 =  x_525 & ~n_16917;
assign n_18301 =  x_1005 & ~n_18254;
assign n_18302 = ~x_1005 &  n_18254;
assign n_18303 =  n_16925 & ~n_18302;
assign n_18304 = ~n_18301 &  n_18303;
assign n_18305 = ~n_18300 & ~n_18304;
assign n_18306 = ~n_18299 &  n_18305;
assign n_18307 = ~x_45 &  n_18259;
assign n_18308 =  x_45 & ~n_18259;
assign n_18309 = ~n_18307 & ~n_18308;
assign n_18310 = ~n_18263 & ~n_18267;
assign n_18311 =  n_18309 & ~n_18310;
assign n_18312 = ~n_18309 &  n_18310;
assign n_18313 = ~n_18311 & ~n_18312;
assign n_18314 = ~x_1933 & ~n_18313;
assign n_18315 =  x_1933 & ~n_18312;
assign n_18316 = ~n_18311 &  n_18315;
assign n_18317 =  n_16920 & ~n_18316;
assign n_18318 = ~n_18314 &  n_18317;
assign n_18319 = ~x_2605 &  n_18271;
assign n_18320 =  x_2605 & ~n_18271;
assign n_18321 = ~n_18319 & ~n_18320;
assign n_18322 = ~n_18275 & ~n_18279;
assign n_18323 =  n_18321 & ~n_18322;
assign n_18324 = ~n_18321 &  n_18322;
assign n_18325 = ~n_18323 & ~n_18324;
assign n_18326 = ~x_2541 & ~n_18325;
assign n_18327 =  x_2541 & ~n_18324;
assign n_18328 = ~n_18323 &  n_18327;
assign n_18329 =  n_16932 & ~n_18328;
assign n_18330 = ~n_18326 &  n_18329;
assign n_18331 = ~n_18318 & ~n_18330;
assign n_18332 =  n_18306 &  n_18331;
assign n_18333 =  x_525 & ~n_18332;
assign n_18334 = ~x_525 &  n_18332;
assign n_18335 = ~n_18333 & ~n_18334;
assign n_18336 = ~x_1644 &  n_18288;
assign n_18337 =  x_1644 & ~n_18288;
assign n_18338 = ~n_18336 & ~n_18337;
assign n_18339 = ~n_18292 & ~n_18296;
assign n_18340 =  n_18338 & ~n_18339;
assign n_18341 = ~n_18338 &  n_18339;
assign n_18342 = ~n_18340 & ~n_18341;
assign n_18343 = ~x_268 & ~n_18342;
assign n_18344 =  x_268 & ~n_18341;
assign n_18345 = ~n_18340 &  n_18344;
assign n_18346 =  n_16927 & ~n_18345;
assign n_18347 = ~n_18343 &  n_18346;
assign n_18348 =  x_524 & ~n_16917;
assign n_18349 =  x_1004 & ~n_18302;
assign n_18350 = ~x_1004 &  n_18302;
assign n_18351 =  n_16925 & ~n_18350;
assign n_18352 = ~n_18349 &  n_18351;
assign n_18353 = ~n_18348 & ~n_18352;
assign n_18354 = ~n_18347 &  n_18353;
assign n_18355 = ~x_44 &  n_18307;
assign n_18356 =  x_44 & ~n_18307;
assign n_18357 = ~n_18355 & ~n_18356;
assign n_18358 = ~n_18311 & ~n_18315;
assign n_18359 =  n_18357 & ~n_18358;
assign n_18360 = ~n_18357 &  n_18358;
assign n_18361 = ~n_18359 & ~n_18360;
assign n_18362 = ~x_1932 & ~n_18361;
assign n_18363 =  x_1932 & ~n_18360;
assign n_18364 = ~n_18359 &  n_18363;
assign n_18365 =  n_16920 & ~n_18364;
assign n_18366 = ~n_18362 &  n_18365;
assign n_18367 = ~x_2604 &  n_18319;
assign n_18368 =  x_2604 & ~n_18319;
assign n_18369 = ~n_18367 & ~n_18368;
assign n_18370 = ~n_18323 & ~n_18327;
assign n_18371 =  n_18369 & ~n_18370;
assign n_18372 = ~n_18369 &  n_18370;
assign n_18373 = ~n_18371 & ~n_18372;
assign n_18374 = ~x_2540 & ~n_18373;
assign n_18375 =  x_2540 & ~n_18372;
assign n_18376 = ~n_18371 &  n_18375;
assign n_18377 =  n_16932 & ~n_18376;
assign n_18378 = ~n_18374 &  n_18377;
assign n_18379 = ~n_18366 & ~n_18378;
assign n_18380 =  n_18354 &  n_18379;
assign n_18381 =  x_524 & ~n_18380;
assign n_18382 = ~x_524 &  n_18380;
assign n_18383 = ~n_18381 & ~n_18382;
assign n_18384 = ~n_18359 & ~n_18363;
assign n_18385 =  x_43 & ~x_1931;
assign n_18386 = ~x_43 &  x_1931;
assign n_18387 = ~n_18385 & ~n_18386;
assign n_18388 =  n_18355 &  n_18387;
assign n_18389 = ~n_18355 & ~n_18387;
assign n_18390 = ~n_18388 & ~n_18389;
assign n_18391 =  n_18384 & ~n_18390;
assign n_18392 = ~n_18384 &  n_18390;
assign n_18393 =  n_16920 & ~n_18392;
assign n_18394 = ~n_18391 &  n_18393;
assign n_18395 =  x_523 & ~n_16917;
assign n_18396 = ~x_1003 &  n_18350;
assign n_18397 =  x_1003 & ~n_18350;
assign n_18398 =  n_16925 & ~n_18397;
assign n_18399 = ~n_18396 &  n_18398;
assign n_18400 = ~n_18395 & ~n_18399;
assign n_18401 = ~n_18394 &  n_18400;
assign n_18402 = ~n_18371 & ~n_18375;
assign n_18403 =  x_2539 & ~x_2603;
assign n_18404 = ~x_2539 &  x_2603;
assign n_18405 = ~n_18403 & ~n_18404;
assign n_18406 =  n_18367 &  n_18405;
assign n_18407 = ~n_18367 & ~n_18405;
assign n_18408 = ~n_18406 & ~n_18407;
assign n_18409 =  n_18402 & ~n_18408;
assign n_18410 = ~n_18402 &  n_18408;
assign n_18411 =  n_16932 & ~n_18410;
assign n_18412 = ~n_18409 &  n_18411;
assign n_18413 = ~n_18340 & ~n_18344;
assign n_18414 =  x_267 & ~x_1643;
assign n_18415 = ~x_267 &  x_1643;
assign n_18416 = ~n_18414 & ~n_18415;
assign n_18417 =  n_18336 &  n_18416;
assign n_18418 = ~n_18336 & ~n_18416;
assign n_18419 = ~n_18417 & ~n_18418;
assign n_18420 =  n_18413 & ~n_18419;
assign n_18421 = ~n_18413 &  n_18419;
assign n_18422 =  n_16927 & ~n_18421;
assign n_18423 = ~n_18420 &  n_18422;
assign n_18424 = ~n_18412 & ~n_18423;
assign n_18425 =  n_18401 &  n_18424;
assign n_18426 =  x_523 & ~n_18425;
assign n_18427 = ~x_523 &  n_18425;
assign n_18428 = ~n_18426 & ~n_18427;
assign n_18429 = ~n_1904 & ~n_13015;
assign n_18430 = ~n_12032 &  n_18429;
assign n_18431 =  n_13012 & ~n_18430;
assign n_18432 =  x_522 & ~n_18431;
assign n_18433 =  x_39 &  n_1904;
assign n_18434 =  n_13012 &  n_18433;
assign n_18435 =  x_138 &  x_2858;
assign n_18436 = ~x_138 & ~x_2858;
assign n_18437 = ~n_18435 & ~n_18436;
assign n_18438 =  n_18434 &  n_18437;
assign n_18439 =  n_2100 &  n_982;
assign n_18440 =  n_12420 &  n_18439;
assign n_18441 =  x_330 &  x_394;
assign n_18442 = ~x_330 & ~x_394;
assign n_18443 = ~n_18441 & ~n_18442;
assign n_18444 =  n_18440 &  n_18443;
assign n_18445 =  n_10319 &  n_13012;
assign n_18446 =  n_1903 &  n_18445;
assign n_18447 =  x_1066 &  n_18446;
assign n_18448 =  n_12420 &  n_1904;
assign n_18449 =  x_650 &  x_2058;
assign n_18450 = ~x_650 & ~x_2058;
assign n_18451 = ~n_18449 & ~n_18450;
assign n_18452 =  n_18448 &  n_18451;
assign n_18453 = ~n_18447 & ~n_18452;
assign n_18454 = ~n_18444 &  n_18453;
assign n_18455 = ~n_18438 &  n_18454;
assign n_18456 = ~n_18432 &  n_18455;
assign n_18457 =  x_522 & ~n_18456;
assign n_18458 = ~x_522 &  n_18456;
assign n_18459 = ~n_18457 & ~n_18458;
assign n_18460 =  x_521 & ~n_18431;
assign n_18461 = ~x_2057 & ~x_2058;
assign n_18462 =  x_2057 &  x_2058;
assign n_18463 = ~n_18461 & ~n_18462;
assign n_18464 =  x_649 &  n_18463;
assign n_18465 = ~x_649 & ~n_18463;
assign n_18466 = ~n_18464 & ~n_18465;
assign n_18467 = ~n_18449 & ~n_18466;
assign n_18468 =  n_18449 &  n_18466;
assign n_18469 =  n_18448 & ~n_18468;
assign n_18470 = ~n_18467 &  n_18469;
assign n_18471 = ~x_1065 & ~x_1066;
assign n_18472 =  x_1065 &  x_1066;
assign n_18473 = ~n_18471 & ~n_18472;
assign n_18474 =  n_18446 &  n_18473;
assign n_18475 = ~n_18470 & ~n_18474;
assign n_18476 = ~x_393 & ~x_394;
assign n_18477 =  x_393 &  x_394;
assign n_18478 = ~n_18476 & ~n_18477;
assign n_18479 =  x_329 &  n_18478;
assign n_18480 = ~x_329 & ~n_18478;
assign n_18481 = ~n_18479 & ~n_18480;
assign n_18482 = ~n_18441 & ~n_18481;
assign n_18483 =  n_18441 &  n_18481;
assign n_18484 =  n_18440 & ~n_18483;
assign n_18485 = ~n_18482 &  n_18484;
assign n_18486 = ~x_137 & ~x_138;
assign n_18487 =  x_137 &  x_138;
assign n_18488 = ~n_18486 & ~n_18487;
assign n_18489 =  x_2857 &  n_18488;
assign n_18490 = ~x_2857 & ~n_18488;
assign n_18491 = ~n_18489 & ~n_18490;
assign n_18492 =  n_18435 &  n_18491;
assign n_18493 = ~n_18435 & ~n_18491;
assign n_18494 = ~n_18492 & ~n_18493;
assign n_18495 =  n_18434 &  n_18494;
assign n_18496 = ~n_18485 & ~n_18495;
assign n_18497 =  n_18475 &  n_18496;
assign n_18498 = ~n_18460 &  n_18497;
assign n_18499 =  x_521 & ~n_18498;
assign n_18500 = ~x_521 &  n_18498;
assign n_18501 = ~n_18499 & ~n_18500;
assign n_18502 = ~x_392 &  n_18476;
assign n_18503 =  x_392 & ~n_18476;
assign n_18504 = ~n_18502 & ~n_18503;
assign n_18505 = ~x_329 &  x_393;
assign n_18506 =  n_18441 & ~n_18505;
assign n_18507 = ~n_18506 & ~n_18479;
assign n_18508 =  n_18504 & ~n_18507;
assign n_18509 = ~n_18504 &  n_18507;
assign n_18510 = ~n_18508 & ~n_18509;
assign n_18511 = ~x_328 & ~n_18510;
assign n_18512 =  x_328 & ~n_18509;
assign n_18513 = ~n_18508 &  n_18512;
assign n_18514 =  n_18440 & ~n_18513;
assign n_18515 = ~n_18511 &  n_18514;
assign n_18516 =  x_520 & ~n_18431;
assign n_18517 = ~x_1064 &  n_18471;
assign n_18518 =  x_1064 & ~n_18471;
assign n_18519 = ~n_18517 & ~n_18518;
assign n_18520 =  n_18446 &  n_18519;
assign n_18521 = ~n_18516 & ~n_18520;
assign n_18522 = ~n_18515 &  n_18521;
assign n_18523 = ~x_2056 &  n_18461;
assign n_18524 =  x_2056 & ~n_18461;
assign n_18525 = ~n_18523 & ~n_18524;
assign n_18526 = ~x_649 &  x_2057;
assign n_18527 =  n_18449 & ~n_18526;
assign n_18528 = ~n_18527 & ~n_18464;
assign n_18529 =  n_18525 & ~n_18528;
assign n_18530 = ~n_18525 &  n_18528;
assign n_18531 = ~n_18529 & ~n_18530;
assign n_18532 = ~x_648 & ~n_18531;
assign n_18533 =  x_648 & ~n_18530;
assign n_18534 = ~n_18529 &  n_18533;
assign n_18535 =  n_18448 & ~n_18534;
assign n_18536 = ~n_18532 &  n_18535;
assign n_18537 = ~x_136 &  n_18486;
assign n_18538 =  x_136 & ~n_18486;
assign n_18539 = ~n_18537 & ~n_18538;
assign n_18540 =  x_137 & ~x_2857;
assign n_18541 =  n_18435 & ~n_18540;
assign n_18542 = ~n_18541 & ~n_18489;
assign n_18543 =  n_18539 & ~n_18542;
assign n_18544 = ~n_18539 &  n_18542;
assign n_18545 = ~n_18543 & ~n_18544;
assign n_18546 = ~x_2856 & ~n_18545;
assign n_18547 =  x_2856 & ~n_18544;
assign n_18548 = ~n_18543 &  n_18547;
assign n_18549 =  n_18434 & ~n_18548;
assign n_18550 = ~n_18546 &  n_18549;
assign n_18551 = ~n_18536 & ~n_18550;
assign n_18552 =  n_18522 &  n_18551;
assign n_18553 =  x_520 & ~n_18552;
assign n_18554 = ~x_520 &  n_18552;
assign n_18555 = ~n_18553 & ~n_18554;
assign n_18556 = ~x_391 &  n_18502;
assign n_18557 =  x_391 & ~n_18502;
assign n_18558 = ~n_18556 & ~n_18557;
assign n_18559 = ~n_18508 & ~n_18512;
assign n_18560 =  n_18558 & ~n_18559;
assign n_18561 = ~n_18558 &  n_18559;
assign n_18562 = ~n_18560 & ~n_18561;
assign n_18563 = ~x_327 & ~n_18562;
assign n_18564 =  x_327 & ~n_18561;
assign n_18565 = ~n_18560 &  n_18564;
assign n_18566 =  n_18440 & ~n_18565;
assign n_18567 = ~n_18563 &  n_18566;
assign n_18568 =  x_519 & ~n_18431;
assign n_18569 = ~x_1063 &  n_18517;
assign n_18570 =  x_1063 & ~n_18517;
assign n_18571 = ~n_18569 & ~n_18570;
assign n_18572 =  n_18446 &  n_18571;
assign n_18573 = ~n_18568 & ~n_18572;
assign n_18574 = ~n_18567 &  n_18573;
assign n_18575 = ~x_135 &  n_18537;
assign n_18576 =  x_135 & ~n_18537;
assign n_18577 = ~n_18575 & ~n_18576;
assign n_18578 = ~n_18543 & ~n_18547;
assign n_18579 =  n_18577 & ~n_18578;
assign n_18580 = ~n_18577 &  n_18578;
assign n_18581 = ~n_18579 & ~n_18580;
assign n_18582 = ~x_2855 & ~n_18581;
assign n_18583 =  x_2855 &  n_18581;
assign n_18584 =  n_18434 & ~n_18583;
assign n_18585 = ~n_18582 &  n_18584;
assign n_18586 = ~x_2055 &  n_18523;
assign n_18587 =  x_2055 & ~n_18523;
assign n_18588 = ~n_18586 & ~n_18587;
assign n_18589 = ~n_18529 & ~n_18533;
assign n_18590 =  n_18588 & ~n_18589;
assign n_18591 = ~n_18588 &  n_18589;
assign n_18592 = ~n_18590 & ~n_18591;
assign n_18593 = ~x_647 & ~n_18592;
assign n_18594 =  x_647 & ~n_18591;
assign n_18595 = ~n_18590 &  n_18594;
assign n_18596 =  n_18448 & ~n_18595;
assign n_18597 = ~n_18593 &  n_18596;
assign n_18598 = ~n_18585 & ~n_18597;
assign n_18599 =  n_18574 &  n_18598;
assign n_18600 =  x_519 & ~n_18599;
assign n_18601 = ~x_519 &  n_18599;
assign n_18602 = ~n_18600 & ~n_18601;
assign n_18603 = ~x_390 &  n_18556;
assign n_18604 =  x_390 & ~n_18556;
assign n_18605 = ~n_18603 & ~n_18604;
assign n_18606 = ~n_18560 & ~n_18564;
assign n_18607 =  n_18605 & ~n_18606;
assign n_18608 = ~n_18605 &  n_18606;
assign n_18609 = ~n_18607 & ~n_18608;
assign n_18610 = ~x_326 & ~n_18609;
assign n_18611 =  x_326 & ~n_18608;
assign n_18612 = ~n_18607 &  n_18611;
assign n_18613 =  n_18440 & ~n_18612;
assign n_18614 = ~n_18610 &  n_18613;
assign n_18615 =  x_518 & ~n_18431;
assign n_18616 =  x_1062 & ~n_18569;
assign n_18617 = ~x_1062 &  n_18569;
assign n_18618 =  n_18446 & ~n_18617;
assign n_18619 = ~n_18616 &  n_18618;
assign n_18620 = ~n_18615 & ~n_18619;
assign n_18621 = ~n_18614 &  n_18620;
assign n_18622 = ~x_134 &  n_18575;
assign n_18623 =  x_134 & ~n_18575;
assign n_18624 = ~n_18622 & ~n_18623;
assign n_18625 =  x_2855 & ~n_18580;
assign n_18626 = ~n_18579 & ~n_18625;
assign n_18627 =  n_18624 & ~n_18626;
assign n_18628 = ~n_18624 &  n_18626;
assign n_18629 = ~n_18627 & ~n_18628;
assign n_18630 = ~x_2854 & ~n_18629;
assign n_18631 =  x_2854 &  n_18629;
assign n_18632 =  n_18434 & ~n_18631;
assign n_18633 = ~n_18630 &  n_18632;
assign n_18634 = ~x_2054 &  n_18586;
assign n_18635 =  x_2054 & ~n_18586;
assign n_18636 = ~n_18634 & ~n_18635;
assign n_18637 = ~n_18590 & ~n_18594;
assign n_18638 =  n_18636 & ~n_18637;
assign n_18639 = ~n_18636 &  n_18637;
assign n_18640 = ~n_18638 & ~n_18639;
assign n_18641 = ~x_646 & ~n_18640;
assign n_18642 =  x_646 & ~n_18639;
assign n_18643 = ~n_18638 &  n_18642;
assign n_18644 =  n_18448 & ~n_18643;
assign n_18645 = ~n_18641 &  n_18644;
assign n_18646 = ~n_18633 & ~n_18645;
assign n_18647 =  n_18621 &  n_18646;
assign n_18648 =  x_518 & ~n_18647;
assign n_18649 = ~x_518 &  n_18647;
assign n_18650 = ~n_18648 & ~n_18649;
assign n_18651 = ~x_389 &  n_18603;
assign n_18652 =  x_389 & ~n_18603;
assign n_18653 = ~n_18651 & ~n_18652;
assign n_18654 = ~n_18607 & ~n_18611;
assign n_18655 =  n_18653 & ~n_18654;
assign n_18656 = ~n_18653 &  n_18654;
assign n_18657 = ~n_18655 & ~n_18656;
assign n_18658 = ~x_325 & ~n_18657;
assign n_18659 =  x_325 & ~n_18656;
assign n_18660 = ~n_18655 &  n_18659;
assign n_18661 =  n_18440 & ~n_18660;
assign n_18662 = ~n_18658 &  n_18661;
assign n_18663 =  x_517 & ~n_18431;
assign n_18664 =  x_1061 & ~n_18617;
assign n_18665 = ~x_1061 &  n_18617;
assign n_18666 =  n_18446 & ~n_18665;
assign n_18667 = ~n_18664 &  n_18666;
assign n_18668 = ~n_18663 & ~n_18667;
assign n_18669 = ~n_18662 &  n_18668;
assign n_18670 = ~x_133 &  n_18622;
assign n_18671 =  x_133 & ~n_18622;
assign n_18672 = ~n_18670 & ~n_18671;
assign n_18673 =  x_2854 & ~n_18628;
assign n_18674 = ~n_18627 & ~n_18673;
assign n_18675 =  n_18672 & ~n_18674;
assign n_18676 = ~n_18672 &  n_18674;
assign n_18677 = ~n_18675 & ~n_18676;
assign n_18678 = ~x_2853 & ~n_18677;
assign n_18679 =  x_2853 &  n_18677;
assign n_18680 =  n_18434 & ~n_18679;
assign n_18681 = ~n_18678 &  n_18680;
assign n_18682 = ~x_2053 &  n_18634;
assign n_18683 =  x_2053 & ~n_18634;
assign n_18684 = ~n_18682 & ~n_18683;
assign n_18685 = ~n_18638 & ~n_18642;
assign n_18686 =  n_18684 & ~n_18685;
assign n_18687 = ~n_18684 &  n_18685;
assign n_18688 = ~n_18686 & ~n_18687;
assign n_18689 = ~x_645 & ~n_18688;
assign n_18690 =  x_645 & ~n_18687;
assign n_18691 = ~n_18686 &  n_18690;
assign n_18692 =  n_18448 & ~n_18691;
assign n_18693 = ~n_18689 &  n_18692;
assign n_18694 = ~n_18681 & ~n_18693;
assign n_18695 =  n_18669 &  n_18694;
assign n_18696 =  x_517 & ~n_18695;
assign n_18697 = ~x_517 &  n_18695;
assign n_18698 = ~n_18696 & ~n_18697;
assign n_18699 = ~x_388 &  n_18651;
assign n_18700 =  x_388 & ~n_18651;
assign n_18701 = ~n_18699 & ~n_18700;
assign n_18702 = ~n_18655 & ~n_18659;
assign n_18703 =  n_18701 & ~n_18702;
assign n_18704 = ~n_18701 &  n_18702;
assign n_18705 = ~n_18703 & ~n_18704;
assign n_18706 = ~x_324 & ~n_18705;
assign n_18707 =  x_324 & ~n_18704;
assign n_18708 = ~n_18703 &  n_18707;
assign n_18709 =  n_18440 & ~n_18708;
assign n_18710 = ~n_18706 &  n_18709;
assign n_18711 =  x_516 & ~n_18431;
assign n_18712 =  x_1060 & ~n_18665;
assign n_18713 = ~x_1060 &  n_18665;
assign n_18714 =  n_18446 & ~n_18713;
assign n_18715 = ~n_18712 &  n_18714;
assign n_18716 = ~n_18711 & ~n_18715;
assign n_18717 = ~n_18710 &  n_18716;
assign n_18718 = ~x_132 &  n_18670;
assign n_18719 =  x_132 & ~n_18670;
assign n_18720 = ~n_18718 & ~n_18719;
assign n_18721 =  x_2853 & ~n_18676;
assign n_18722 = ~n_18675 & ~n_18721;
assign n_18723 =  n_18720 & ~n_18722;
assign n_18724 = ~n_18720 &  n_18722;
assign n_18725 = ~n_18723 & ~n_18724;
assign n_18726 = ~x_2852 & ~n_18725;
assign n_18727 =  x_2852 &  n_18725;
assign n_18728 =  n_18434 & ~n_18727;
assign n_18729 = ~n_18726 &  n_18728;
assign n_18730 = ~x_2052 &  n_18682;
assign n_18731 =  x_2052 & ~n_18682;
assign n_18732 = ~n_18730 & ~n_18731;
assign n_18733 = ~n_18686 & ~n_18690;
assign n_18734 =  n_18732 & ~n_18733;
assign n_18735 = ~n_18732 &  n_18733;
assign n_18736 = ~n_18734 & ~n_18735;
assign n_18737 = ~x_644 & ~n_18736;
assign n_18738 =  x_644 & ~n_18735;
assign n_18739 = ~n_18734 &  n_18738;
assign n_18740 =  n_18448 & ~n_18739;
assign n_18741 = ~n_18737 &  n_18740;
assign n_18742 = ~n_18729 & ~n_18741;
assign n_18743 =  n_18717 &  n_18742;
assign n_18744 =  x_516 & ~n_18743;
assign n_18745 = ~x_516 &  n_18743;
assign n_18746 = ~n_18744 & ~n_18745;
assign n_18747 = ~x_387 &  n_18699;
assign n_18748 =  x_387 & ~n_18699;
assign n_18749 = ~n_18747 & ~n_18748;
assign n_18750 = ~n_18703 & ~n_18707;
assign n_18751 =  n_18749 & ~n_18750;
assign n_18752 = ~n_18749 &  n_18750;
assign n_18753 = ~n_18751 & ~n_18752;
assign n_18754 = ~x_323 & ~n_18753;
assign n_18755 =  x_323 & ~n_18752;
assign n_18756 = ~n_18751 &  n_18755;
assign n_18757 =  n_18440 & ~n_18756;
assign n_18758 = ~n_18754 &  n_18757;
assign n_18759 =  x_515 & ~n_18431;
assign n_18760 =  x_1059 & ~n_18713;
assign n_18761 = ~x_1059 &  n_18713;
assign n_18762 =  n_18446 & ~n_18761;
assign n_18763 = ~n_18760 &  n_18762;
assign n_18764 = ~n_18759 & ~n_18763;
assign n_18765 = ~n_18758 &  n_18764;
assign n_18766 = ~x_131 &  n_18718;
assign n_18767 =  x_131 & ~n_18718;
assign n_18768 = ~n_18766 & ~n_18767;
assign n_18769 =  x_2852 & ~n_18724;
assign n_18770 = ~n_18723 & ~n_18769;
assign n_18771 =  n_18768 & ~n_18770;
assign n_18772 = ~n_18768 &  n_18770;
assign n_18773 = ~n_18771 & ~n_18772;
assign n_18774 = ~x_2851 & ~n_18773;
assign n_18775 =  x_2851 &  n_18773;
assign n_18776 =  n_18434 & ~n_18775;
assign n_18777 = ~n_18774 &  n_18776;
assign n_18778 = ~x_2051 &  n_18730;
assign n_18779 =  x_2051 & ~n_18730;
assign n_18780 = ~n_18778 & ~n_18779;
assign n_18781 = ~n_18734 & ~n_18738;
assign n_18782 =  n_18780 & ~n_18781;
assign n_18783 = ~n_18780 &  n_18781;
assign n_18784 = ~n_18782 & ~n_18783;
assign n_18785 = ~x_643 & ~n_18784;
assign n_18786 =  x_643 & ~n_18783;
assign n_18787 = ~n_18782 &  n_18786;
assign n_18788 =  n_18448 & ~n_18787;
assign n_18789 = ~n_18785 &  n_18788;
assign n_18790 = ~n_18777 & ~n_18789;
assign n_18791 =  n_18765 &  n_18790;
assign n_18792 =  x_515 & ~n_18791;
assign n_18793 = ~x_515 &  n_18791;
assign n_18794 = ~n_18792 & ~n_18793;
assign n_18795 = ~x_386 &  n_18747;
assign n_18796 =  x_386 & ~n_18747;
assign n_18797 = ~n_18795 & ~n_18796;
assign n_18798 = ~n_18751 & ~n_18755;
assign n_18799 =  n_18797 & ~n_18798;
assign n_18800 = ~n_18797 &  n_18798;
assign n_18801 = ~n_18799 & ~n_18800;
assign n_18802 = ~x_322 & ~n_18801;
assign n_18803 =  x_322 & ~n_18800;
assign n_18804 = ~n_18799 &  n_18803;
assign n_18805 =  n_18440 & ~n_18804;
assign n_18806 = ~n_18802 &  n_18805;
assign n_18807 =  x_514 & ~n_18431;
assign n_18808 =  x_1058 & ~n_18761;
assign n_18809 = ~x_1058 &  n_18761;
assign n_18810 =  n_18446 & ~n_18809;
assign n_18811 = ~n_18808 &  n_18810;
assign n_18812 = ~n_18807 & ~n_18811;
assign n_18813 = ~n_18806 &  n_18812;
assign n_18814 = ~x_130 &  n_18766;
assign n_18815 =  x_130 & ~n_18766;
assign n_18816 = ~n_18814 & ~n_18815;
assign n_18817 =  x_2851 & ~n_18772;
assign n_18818 = ~n_18771 & ~n_18817;
assign n_18819 =  n_18816 & ~n_18818;
assign n_18820 = ~n_18816 &  n_18818;
assign n_18821 = ~n_18819 & ~n_18820;
assign n_18822 = ~x_2850 & ~n_18821;
assign n_18823 =  x_2850 &  n_18821;
assign n_18824 =  n_18434 & ~n_18823;
assign n_18825 = ~n_18822 &  n_18824;
assign n_18826 = ~x_2050 &  n_18778;
assign n_18827 =  x_2050 & ~n_18778;
assign n_18828 = ~n_18826 & ~n_18827;
assign n_18829 = ~n_18782 & ~n_18786;
assign n_18830 =  n_18828 & ~n_18829;
assign n_18831 = ~n_18828 &  n_18829;
assign n_18832 = ~n_18830 & ~n_18831;
assign n_18833 = ~x_642 & ~n_18832;
assign n_18834 =  x_642 & ~n_18831;
assign n_18835 = ~n_18830 &  n_18834;
assign n_18836 =  n_18448 & ~n_18835;
assign n_18837 = ~n_18833 &  n_18836;
assign n_18838 = ~n_18825 & ~n_18837;
assign n_18839 =  n_18813 &  n_18838;
assign n_18840 =  x_514 & ~n_18839;
assign n_18841 = ~x_514 &  n_18839;
assign n_18842 = ~n_18840 & ~n_18841;
assign n_18843 = ~x_385 &  n_18795;
assign n_18844 =  x_385 & ~n_18795;
assign n_18845 = ~n_18843 & ~n_18844;
assign n_18846 = ~n_18799 & ~n_18803;
assign n_18847 =  n_18845 & ~n_18846;
assign n_18848 = ~n_18845 &  n_18846;
assign n_18849 = ~n_18847 & ~n_18848;
assign n_18850 = ~x_321 & ~n_18849;
assign n_18851 =  x_321 & ~n_18848;
assign n_18852 = ~n_18847 &  n_18851;
assign n_18853 =  n_18440 & ~n_18852;
assign n_18854 = ~n_18850 &  n_18853;
assign n_18855 =  x_513 & ~n_18431;
assign n_18856 =  x_1057 & ~n_18809;
assign n_18857 = ~x_1057 &  n_18809;
assign n_18858 =  n_18446 & ~n_18857;
assign n_18859 = ~n_18856 &  n_18858;
assign n_18860 = ~n_18855 & ~n_18859;
assign n_18861 = ~n_18854 &  n_18860;
assign n_18862 = ~x_129 &  n_18814;
assign n_18863 =  x_129 & ~n_18814;
assign n_18864 = ~n_18862 & ~n_18863;
assign n_18865 =  x_2850 & ~n_18820;
assign n_18866 = ~n_18819 & ~n_18865;
assign n_18867 =  n_18864 & ~n_18866;
assign n_18868 = ~n_18864 &  n_18866;
assign n_18869 = ~n_18867 & ~n_18868;
assign n_18870 = ~x_2849 & ~n_18869;
assign n_18871 =  x_2849 &  n_18869;
assign n_18872 =  n_18434 & ~n_18871;
assign n_18873 = ~n_18870 &  n_18872;
assign n_18874 = ~x_2049 &  n_18826;
assign n_18875 =  x_2049 & ~n_18826;
assign n_18876 = ~n_18874 & ~n_18875;
assign n_18877 = ~n_18830 & ~n_18834;
assign n_18878 =  n_18876 & ~n_18877;
assign n_18879 = ~n_18876 &  n_18877;
assign n_18880 = ~n_18878 & ~n_18879;
assign n_18881 = ~x_641 & ~n_18880;
assign n_18882 =  x_641 & ~n_18879;
assign n_18883 = ~n_18878 &  n_18882;
assign n_18884 =  n_18448 & ~n_18883;
assign n_18885 = ~n_18881 &  n_18884;
assign n_18886 = ~n_18873 & ~n_18885;
assign n_18887 =  n_18861 &  n_18886;
assign n_18888 =  x_513 & ~n_18887;
assign n_18889 = ~x_513 &  n_18887;
assign n_18890 = ~n_18888 & ~n_18889;
assign n_18891 = ~x_384 &  n_18843;
assign n_18892 =  x_384 & ~n_18843;
assign n_18893 = ~n_18891 & ~n_18892;
assign n_18894 = ~n_18847 & ~n_18851;
assign n_18895 =  n_18893 & ~n_18894;
assign n_18896 = ~n_18893 &  n_18894;
assign n_18897 = ~n_18895 & ~n_18896;
assign n_18898 = ~x_320 & ~n_18897;
assign n_18899 =  x_320 & ~n_18896;
assign n_18900 = ~n_18895 &  n_18899;
assign n_18901 =  n_18440 & ~n_18900;
assign n_18902 = ~n_18898 &  n_18901;
assign n_18903 =  x_512 & ~n_18431;
assign n_18904 =  x_1056 & ~n_18857;
assign n_18905 = ~x_1056 &  n_18857;
assign n_18906 =  n_18446 & ~n_18905;
assign n_18907 = ~n_18904 &  n_18906;
assign n_18908 = ~n_18903 & ~n_18907;
assign n_18909 = ~n_18902 &  n_18908;
assign n_18910 = ~x_128 &  n_18862;
assign n_18911 =  x_128 & ~n_18862;
assign n_18912 = ~n_18910 & ~n_18911;
assign n_18913 =  x_2849 & ~n_18868;
assign n_18914 = ~n_18867 & ~n_18913;
assign n_18915 =  n_18912 & ~n_18914;
assign n_18916 = ~n_18912 &  n_18914;
assign n_18917 = ~n_18915 & ~n_18916;
assign n_18918 = ~x_2848 & ~n_18917;
assign n_18919 =  x_2848 &  n_18917;
assign n_18920 =  n_18434 & ~n_18919;
assign n_18921 = ~n_18918 &  n_18920;
assign n_18922 = ~x_2048 &  n_18874;
assign n_18923 =  x_2048 & ~n_18874;
assign n_18924 = ~n_18922 & ~n_18923;
assign n_18925 = ~n_18878 & ~n_18882;
assign n_18926 =  n_18924 & ~n_18925;
assign n_18927 = ~n_18924 &  n_18925;
assign n_18928 = ~n_18926 & ~n_18927;
assign n_18929 = ~x_640 & ~n_18928;
assign n_18930 =  x_640 & ~n_18927;
assign n_18931 = ~n_18926 &  n_18930;
assign n_18932 =  n_18448 & ~n_18931;
assign n_18933 = ~n_18929 &  n_18932;
assign n_18934 = ~n_18921 & ~n_18933;
assign n_18935 =  n_18909 &  n_18934;
assign n_18936 =  x_512 & ~n_18935;
assign n_18937 = ~x_512 &  n_18935;
assign n_18938 = ~n_18936 & ~n_18937;
assign n_18939 = ~x_383 &  n_18891;
assign n_18940 =  x_383 & ~n_18891;
assign n_18941 = ~n_18939 & ~n_18940;
assign n_18942 = ~n_18895 & ~n_18899;
assign n_18943 =  n_18941 & ~n_18942;
assign n_18944 = ~n_18941 &  n_18942;
assign n_18945 = ~n_18943 & ~n_18944;
assign n_18946 = ~x_319 & ~n_18945;
assign n_18947 =  x_319 & ~n_18944;
assign n_18948 = ~n_18943 &  n_18947;
assign n_18949 =  n_18440 & ~n_18948;
assign n_18950 = ~n_18946 &  n_18949;
assign n_18951 =  x_511 & ~n_18431;
assign n_18952 =  x_1055 & ~n_18905;
assign n_18953 = ~x_1055 &  n_18905;
assign n_18954 =  n_18446 & ~n_18953;
assign n_18955 = ~n_18952 &  n_18954;
assign n_18956 = ~n_18951 & ~n_18955;
assign n_18957 = ~n_18950 &  n_18956;
assign n_18958 = ~x_127 &  n_18910;
assign n_18959 =  x_127 & ~n_18910;
assign n_18960 = ~n_18958 & ~n_18959;
assign n_18961 =  x_2848 & ~n_18916;
assign n_18962 = ~n_18915 & ~n_18961;
assign n_18963 =  n_18960 & ~n_18962;
assign n_18964 = ~n_18960 &  n_18962;
assign n_18965 = ~n_18963 & ~n_18964;
assign n_18966 = ~x_2847 & ~n_18965;
assign n_18967 =  x_2847 &  n_18965;
assign n_18968 =  n_18434 & ~n_18967;
assign n_18969 = ~n_18966 &  n_18968;
assign n_18970 = ~x_2047 &  n_18922;
assign n_18971 =  x_2047 & ~n_18922;
assign n_18972 = ~n_18970 & ~n_18971;
assign n_18973 = ~n_18926 & ~n_18930;
assign n_18974 =  n_18972 & ~n_18973;
assign n_18975 = ~n_18972 &  n_18973;
assign n_18976 = ~n_18974 & ~n_18975;
assign n_18977 = ~x_639 & ~n_18976;
assign n_18978 =  x_639 & ~n_18975;
assign n_18979 = ~n_18974 &  n_18978;
assign n_18980 =  n_18448 & ~n_18979;
assign n_18981 = ~n_18977 &  n_18980;
assign n_18982 = ~n_18969 & ~n_18981;
assign n_18983 =  n_18957 &  n_18982;
assign n_18984 =  x_511 & ~n_18983;
assign n_18985 = ~x_511 &  n_18983;
assign n_18986 = ~n_18984 & ~n_18985;
assign n_18987 = ~x_382 &  n_18939;
assign n_18988 =  x_382 & ~n_18939;
assign n_18989 = ~n_18987 & ~n_18988;
assign n_18990 = ~n_18943 & ~n_18947;
assign n_18991 =  n_18989 & ~n_18990;
assign n_18992 = ~n_18989 &  n_18990;
assign n_18993 = ~n_18991 & ~n_18992;
assign n_18994 = ~x_318 & ~n_18993;
assign n_18995 =  x_318 & ~n_18992;
assign n_18996 = ~n_18991 &  n_18995;
assign n_18997 =  n_18440 & ~n_18996;
assign n_18998 = ~n_18994 &  n_18997;
assign n_18999 =  x_510 & ~n_18431;
assign n_19000 =  x_1054 & ~n_18953;
assign n_19001 = ~x_1054 &  n_18953;
assign n_19002 =  n_18446 & ~n_19001;
assign n_19003 = ~n_19000 &  n_19002;
assign n_19004 = ~n_18999 & ~n_19003;
assign n_19005 = ~n_18998 &  n_19004;
assign n_19006 = ~x_126 &  n_18958;
assign n_19007 =  x_126 & ~n_18958;
assign n_19008 = ~n_19006 & ~n_19007;
assign n_19009 =  x_2847 & ~n_18964;
assign n_19010 = ~n_18963 & ~n_19009;
assign n_19011 =  n_19008 & ~n_19010;
assign n_19012 = ~n_19008 &  n_19010;
assign n_19013 = ~n_19011 & ~n_19012;
assign n_19014 = ~x_2846 & ~n_19013;
assign n_19015 =  x_2846 &  n_19013;
assign n_19016 =  n_18434 & ~n_19015;
assign n_19017 = ~n_19014 &  n_19016;
assign n_19018 = ~x_2046 &  n_18970;
assign n_19019 =  x_2046 & ~n_18970;
assign n_19020 = ~n_19018 & ~n_19019;
assign n_19021 = ~n_18974 & ~n_18978;
assign n_19022 =  n_19020 & ~n_19021;
assign n_19023 = ~n_19020 &  n_19021;
assign n_19024 = ~n_19022 & ~n_19023;
assign n_19025 = ~x_638 & ~n_19024;
assign n_19026 =  x_638 & ~n_19023;
assign n_19027 = ~n_19022 &  n_19026;
assign n_19028 =  n_18448 & ~n_19027;
assign n_19029 = ~n_19025 &  n_19028;
assign n_19030 = ~n_19017 & ~n_19029;
assign n_19031 =  n_19005 &  n_19030;
assign n_19032 =  x_510 & ~n_19031;
assign n_19033 = ~x_510 &  n_19031;
assign n_19034 = ~n_19032 & ~n_19033;
assign n_19035 = ~x_381 &  n_18987;
assign n_19036 =  x_381 & ~n_18987;
assign n_19037 = ~n_19035 & ~n_19036;
assign n_19038 = ~n_18991 & ~n_18995;
assign n_19039 =  n_19037 & ~n_19038;
assign n_19040 = ~n_19037 &  n_19038;
assign n_19041 = ~n_19039 & ~n_19040;
assign n_19042 = ~x_317 & ~n_19041;
assign n_19043 =  x_317 & ~n_19040;
assign n_19044 = ~n_19039 &  n_19043;
assign n_19045 =  n_18440 & ~n_19044;
assign n_19046 = ~n_19042 &  n_19045;
assign n_19047 =  x_509 & ~n_18431;
assign n_19048 =  x_1053 & ~n_19001;
assign n_19049 = ~x_1053 &  n_19001;
assign n_19050 =  n_18446 & ~n_19049;
assign n_19051 = ~n_19048 &  n_19050;
assign n_19052 = ~n_19047 & ~n_19051;
assign n_19053 = ~n_19046 &  n_19052;
assign n_19054 = ~x_125 &  n_19006;
assign n_19055 =  x_125 & ~n_19006;
assign n_19056 = ~n_19054 & ~n_19055;
assign n_19057 =  x_2846 & ~n_19012;
assign n_19058 = ~n_19011 & ~n_19057;
assign n_19059 =  n_19056 & ~n_19058;
assign n_19060 = ~n_19056 &  n_19058;
assign n_19061 = ~n_19059 & ~n_19060;
assign n_19062 = ~x_2845 & ~n_19061;
assign n_19063 =  x_2845 &  n_19061;
assign n_19064 =  n_18434 & ~n_19063;
assign n_19065 = ~n_19062 &  n_19064;
assign n_19066 = ~x_2045 &  n_19018;
assign n_19067 =  x_2045 & ~n_19018;
assign n_19068 = ~n_19066 & ~n_19067;
assign n_19069 = ~n_19022 & ~n_19026;
assign n_19070 =  n_19068 & ~n_19069;
assign n_19071 = ~n_19068 &  n_19069;
assign n_19072 = ~n_19070 & ~n_19071;
assign n_19073 = ~x_637 & ~n_19072;
assign n_19074 =  x_637 & ~n_19071;
assign n_19075 = ~n_19070 &  n_19074;
assign n_19076 =  n_18448 & ~n_19075;
assign n_19077 = ~n_19073 &  n_19076;
assign n_19078 = ~n_19065 & ~n_19077;
assign n_19079 =  n_19053 &  n_19078;
assign n_19080 =  x_509 & ~n_19079;
assign n_19081 = ~x_509 &  n_19079;
assign n_19082 = ~n_19080 & ~n_19081;
assign n_19083 = ~x_380 &  n_19035;
assign n_19084 =  x_380 & ~n_19035;
assign n_19085 = ~n_19083 & ~n_19084;
assign n_19086 = ~n_19039 & ~n_19043;
assign n_19087 =  n_19085 & ~n_19086;
assign n_19088 = ~n_19085 &  n_19086;
assign n_19089 = ~n_19087 & ~n_19088;
assign n_19090 = ~x_316 & ~n_19089;
assign n_19091 =  x_316 & ~n_19088;
assign n_19092 = ~n_19087 &  n_19091;
assign n_19093 =  n_18440 & ~n_19092;
assign n_19094 = ~n_19090 &  n_19093;
assign n_19095 =  x_508 & ~n_18431;
assign n_19096 =  x_1052 & ~n_19049;
assign n_19097 = ~x_1052 &  n_19049;
assign n_19098 =  n_18446 & ~n_19097;
assign n_19099 = ~n_19096 &  n_19098;
assign n_19100 = ~n_19095 & ~n_19099;
assign n_19101 = ~n_19094 &  n_19100;
assign n_19102 = ~x_124 &  n_19054;
assign n_19103 =  x_124 & ~n_19054;
assign n_19104 = ~n_19102 & ~n_19103;
assign n_19105 =  x_2845 & ~n_19060;
assign n_19106 = ~n_19059 & ~n_19105;
assign n_19107 =  n_19104 & ~n_19106;
assign n_19108 = ~n_19104 &  n_19106;
assign n_19109 = ~n_19107 & ~n_19108;
assign n_19110 = ~x_2844 & ~n_19109;
assign n_19111 =  x_2844 &  n_19109;
assign n_19112 =  n_18434 & ~n_19111;
assign n_19113 = ~n_19110 &  n_19112;
assign n_19114 = ~x_2044 &  n_19066;
assign n_19115 =  x_2044 & ~n_19066;
assign n_19116 = ~n_19114 & ~n_19115;
assign n_19117 = ~n_19070 & ~n_19074;
assign n_19118 =  n_19116 & ~n_19117;
assign n_19119 = ~n_19116 &  n_19117;
assign n_19120 = ~n_19118 & ~n_19119;
assign n_19121 = ~x_636 & ~n_19120;
assign n_19122 =  x_636 & ~n_19119;
assign n_19123 = ~n_19118 &  n_19122;
assign n_19124 =  n_18448 & ~n_19123;
assign n_19125 = ~n_19121 &  n_19124;
assign n_19126 = ~n_19113 & ~n_19125;
assign n_19127 =  n_19101 &  n_19126;
assign n_19128 =  x_508 & ~n_19127;
assign n_19129 = ~x_508 &  n_19127;
assign n_19130 = ~n_19128 & ~n_19129;
assign n_19131 = ~x_379 &  n_19083;
assign n_19132 =  x_379 & ~n_19083;
assign n_19133 = ~n_19131 & ~n_19132;
assign n_19134 = ~n_19087 & ~n_19091;
assign n_19135 =  n_19133 & ~n_19134;
assign n_19136 = ~n_19133 &  n_19134;
assign n_19137 = ~n_19135 & ~n_19136;
assign n_19138 = ~x_315 & ~n_19137;
assign n_19139 =  x_315 & ~n_19136;
assign n_19140 = ~n_19135 &  n_19139;
assign n_19141 =  n_18440 & ~n_19140;
assign n_19142 = ~n_19138 &  n_19141;
assign n_19143 =  x_507 & ~n_18431;
assign n_19144 =  x_1051 & ~n_19097;
assign n_19145 = ~x_1051 &  n_19097;
assign n_19146 =  n_18446 & ~n_19145;
assign n_19147 = ~n_19144 &  n_19146;
assign n_19148 = ~n_19143 & ~n_19147;
assign n_19149 = ~n_19142 &  n_19148;
assign n_19150 = ~x_123 &  n_19102;
assign n_19151 =  x_123 & ~n_19102;
assign n_19152 = ~n_19150 & ~n_19151;
assign n_19153 =  x_2844 & ~n_19108;
assign n_19154 = ~n_19107 & ~n_19153;
assign n_19155 =  n_19152 & ~n_19154;
assign n_19156 = ~n_19152 &  n_19154;
assign n_19157 = ~n_19155 & ~n_19156;
assign n_19158 = ~x_2843 & ~n_19157;
assign n_19159 =  x_2843 &  n_19157;
assign n_19160 =  n_18434 & ~n_19159;
assign n_19161 = ~n_19158 &  n_19160;
assign n_19162 = ~x_2043 &  n_19114;
assign n_19163 =  x_2043 & ~n_19114;
assign n_19164 = ~n_19162 & ~n_19163;
assign n_19165 = ~n_19118 & ~n_19122;
assign n_19166 =  n_19164 & ~n_19165;
assign n_19167 = ~n_19164 &  n_19165;
assign n_19168 = ~n_19166 & ~n_19167;
assign n_19169 = ~x_635 & ~n_19168;
assign n_19170 =  x_635 & ~n_19167;
assign n_19171 = ~n_19166 &  n_19170;
assign n_19172 =  n_18448 & ~n_19171;
assign n_19173 = ~n_19169 &  n_19172;
assign n_19174 = ~n_19161 & ~n_19173;
assign n_19175 =  n_19149 &  n_19174;
assign n_19176 =  x_507 & ~n_19175;
assign n_19177 = ~x_507 &  n_19175;
assign n_19178 = ~n_19176 & ~n_19177;
assign n_19179 = ~x_378 &  n_19131;
assign n_19180 =  x_378 & ~n_19131;
assign n_19181 = ~n_19179 & ~n_19180;
assign n_19182 = ~n_19135 & ~n_19139;
assign n_19183 =  n_19181 & ~n_19182;
assign n_19184 = ~n_19181 &  n_19182;
assign n_19185 = ~n_19183 & ~n_19184;
assign n_19186 = ~x_314 & ~n_19185;
assign n_19187 =  x_314 & ~n_19184;
assign n_19188 = ~n_19183 &  n_19187;
assign n_19189 =  n_18440 & ~n_19188;
assign n_19190 = ~n_19186 &  n_19189;
assign n_19191 =  x_506 & ~n_18431;
assign n_19192 =  x_1050 & ~n_19145;
assign n_19193 = ~x_1050 &  n_19145;
assign n_19194 =  n_18446 & ~n_19193;
assign n_19195 = ~n_19192 &  n_19194;
assign n_19196 = ~n_19191 & ~n_19195;
assign n_19197 = ~n_19190 &  n_19196;
assign n_19198 = ~x_122 &  n_19150;
assign n_19199 =  x_122 & ~n_19150;
assign n_19200 = ~n_19198 & ~n_19199;
assign n_19201 =  x_2843 & ~n_19156;
assign n_19202 = ~n_19155 & ~n_19201;
assign n_19203 =  n_19200 & ~n_19202;
assign n_19204 = ~n_19200 &  n_19202;
assign n_19205 = ~n_19203 & ~n_19204;
assign n_19206 = ~x_2842 & ~n_19205;
assign n_19207 =  x_2842 &  n_19205;
assign n_19208 =  n_18434 & ~n_19207;
assign n_19209 = ~n_19206 &  n_19208;
assign n_19210 = ~x_2042 &  n_19162;
assign n_19211 =  x_2042 & ~n_19162;
assign n_19212 = ~n_19210 & ~n_19211;
assign n_19213 = ~n_19166 & ~n_19170;
assign n_19214 =  n_19212 & ~n_19213;
assign n_19215 = ~n_19212 &  n_19213;
assign n_19216 = ~n_19214 & ~n_19215;
assign n_19217 = ~x_634 & ~n_19216;
assign n_19218 =  x_634 & ~n_19215;
assign n_19219 = ~n_19214 &  n_19218;
assign n_19220 =  n_18448 & ~n_19219;
assign n_19221 = ~n_19217 &  n_19220;
assign n_19222 = ~n_19209 & ~n_19221;
assign n_19223 =  n_19197 &  n_19222;
assign n_19224 =  x_506 & ~n_19223;
assign n_19225 = ~x_506 &  n_19223;
assign n_19226 = ~n_19224 & ~n_19225;
assign n_19227 = ~x_377 &  n_19179;
assign n_19228 =  x_377 & ~n_19179;
assign n_19229 = ~n_19227 & ~n_19228;
assign n_19230 = ~n_19183 & ~n_19187;
assign n_19231 =  n_19229 & ~n_19230;
assign n_19232 = ~n_19229 &  n_19230;
assign n_19233 = ~n_19231 & ~n_19232;
assign n_19234 = ~x_313 & ~n_19233;
assign n_19235 =  x_313 & ~n_19232;
assign n_19236 = ~n_19231 &  n_19235;
assign n_19237 =  n_18440 & ~n_19236;
assign n_19238 = ~n_19234 &  n_19237;
assign n_19239 =  x_505 & ~n_18431;
assign n_19240 =  x_1049 & ~n_19193;
assign n_19241 = ~x_1049 &  n_19193;
assign n_19242 =  n_18446 & ~n_19241;
assign n_19243 = ~n_19240 &  n_19242;
assign n_19244 = ~n_19239 & ~n_19243;
assign n_19245 = ~n_19238 &  n_19244;
assign n_19246 = ~x_121 &  n_19198;
assign n_19247 =  x_121 & ~n_19198;
assign n_19248 = ~n_19246 & ~n_19247;
assign n_19249 =  x_2842 & ~n_19204;
assign n_19250 = ~n_19203 & ~n_19249;
assign n_19251 =  n_19248 & ~n_19250;
assign n_19252 = ~n_19248 &  n_19250;
assign n_19253 = ~n_19251 & ~n_19252;
assign n_19254 = ~x_2841 & ~n_19253;
assign n_19255 =  x_2841 &  n_19253;
assign n_19256 =  n_18434 & ~n_19255;
assign n_19257 = ~n_19254 &  n_19256;
assign n_19258 = ~x_2041 &  n_19210;
assign n_19259 =  x_2041 & ~n_19210;
assign n_19260 = ~n_19258 & ~n_19259;
assign n_19261 = ~n_19214 & ~n_19218;
assign n_19262 =  n_19260 & ~n_19261;
assign n_19263 = ~n_19260 &  n_19261;
assign n_19264 = ~n_19262 & ~n_19263;
assign n_19265 = ~x_633 & ~n_19264;
assign n_19266 =  x_633 & ~n_19263;
assign n_19267 = ~n_19262 &  n_19266;
assign n_19268 =  n_18448 & ~n_19267;
assign n_19269 = ~n_19265 &  n_19268;
assign n_19270 = ~n_19257 & ~n_19269;
assign n_19271 =  n_19245 &  n_19270;
assign n_19272 =  x_505 & ~n_19271;
assign n_19273 = ~x_505 &  n_19271;
assign n_19274 = ~n_19272 & ~n_19273;
assign n_19275 = ~x_376 &  n_19227;
assign n_19276 =  x_376 & ~n_19227;
assign n_19277 = ~n_19275 & ~n_19276;
assign n_19278 = ~n_19231 & ~n_19235;
assign n_19279 =  n_19277 & ~n_19278;
assign n_19280 = ~n_19277 &  n_19278;
assign n_19281 = ~n_19279 & ~n_19280;
assign n_19282 = ~x_312 & ~n_19281;
assign n_19283 =  x_312 & ~n_19280;
assign n_19284 = ~n_19279 &  n_19283;
assign n_19285 =  n_18440 & ~n_19284;
assign n_19286 = ~n_19282 &  n_19285;
assign n_19287 =  x_504 & ~n_18431;
assign n_19288 =  x_1048 & ~n_19241;
assign n_19289 = ~x_1048 &  n_19241;
assign n_19290 =  n_18446 & ~n_19289;
assign n_19291 = ~n_19288 &  n_19290;
assign n_19292 = ~n_19287 & ~n_19291;
assign n_19293 = ~n_19286 &  n_19292;
assign n_19294 = ~x_120 &  n_19246;
assign n_19295 =  x_120 & ~n_19246;
assign n_19296 = ~n_19294 & ~n_19295;
assign n_19297 =  x_2841 & ~n_19252;
assign n_19298 = ~n_19251 & ~n_19297;
assign n_19299 =  n_19296 & ~n_19298;
assign n_19300 = ~n_19296 &  n_19298;
assign n_19301 = ~n_19299 & ~n_19300;
assign n_19302 = ~x_2840 & ~n_19301;
assign n_19303 =  x_2840 &  n_19301;
assign n_19304 =  n_18434 & ~n_19303;
assign n_19305 = ~n_19302 &  n_19304;
assign n_19306 = ~x_2040 &  n_19258;
assign n_19307 =  x_2040 & ~n_19258;
assign n_19308 = ~n_19306 & ~n_19307;
assign n_19309 = ~n_19262 & ~n_19266;
assign n_19310 =  n_19308 & ~n_19309;
assign n_19311 = ~n_19308 &  n_19309;
assign n_19312 = ~n_19310 & ~n_19311;
assign n_19313 = ~x_632 & ~n_19312;
assign n_19314 =  x_632 & ~n_19311;
assign n_19315 = ~n_19310 &  n_19314;
assign n_19316 =  n_18448 & ~n_19315;
assign n_19317 = ~n_19313 &  n_19316;
assign n_19318 = ~n_19305 & ~n_19317;
assign n_19319 =  n_19293 &  n_19318;
assign n_19320 =  x_504 & ~n_19319;
assign n_19321 = ~x_504 &  n_19319;
assign n_19322 = ~n_19320 & ~n_19321;
assign n_19323 = ~x_375 &  n_19275;
assign n_19324 =  x_375 & ~n_19275;
assign n_19325 = ~n_19323 & ~n_19324;
assign n_19326 = ~n_19279 & ~n_19283;
assign n_19327 =  n_19325 & ~n_19326;
assign n_19328 = ~n_19325 &  n_19326;
assign n_19329 = ~n_19327 & ~n_19328;
assign n_19330 = ~x_311 & ~n_19329;
assign n_19331 =  x_311 & ~n_19328;
assign n_19332 = ~n_19327 &  n_19331;
assign n_19333 =  n_18440 & ~n_19332;
assign n_19334 = ~n_19330 &  n_19333;
assign n_19335 =  x_503 & ~n_18431;
assign n_19336 =  x_1047 & ~n_19289;
assign n_19337 = ~x_1047 &  n_19289;
assign n_19338 =  n_18446 & ~n_19337;
assign n_19339 = ~n_19336 &  n_19338;
assign n_19340 = ~n_19335 & ~n_19339;
assign n_19341 = ~n_19334 &  n_19340;
assign n_19342 = ~x_119 &  n_19294;
assign n_19343 =  x_119 & ~n_19294;
assign n_19344 = ~n_19342 & ~n_19343;
assign n_19345 =  x_2840 & ~n_19300;
assign n_19346 = ~n_19299 & ~n_19345;
assign n_19347 =  n_19344 & ~n_19346;
assign n_19348 = ~n_19344 &  n_19346;
assign n_19349 = ~n_19347 & ~n_19348;
assign n_19350 = ~x_2839 & ~n_19349;
assign n_19351 =  x_2839 &  n_19349;
assign n_19352 =  n_18434 & ~n_19351;
assign n_19353 = ~n_19350 &  n_19352;
assign n_19354 = ~x_2039 &  n_19306;
assign n_19355 =  x_2039 & ~n_19306;
assign n_19356 = ~n_19354 & ~n_19355;
assign n_19357 = ~n_19310 & ~n_19314;
assign n_19358 =  n_19356 & ~n_19357;
assign n_19359 = ~n_19356 &  n_19357;
assign n_19360 = ~n_19358 & ~n_19359;
assign n_19361 = ~x_631 & ~n_19360;
assign n_19362 =  x_631 & ~n_19359;
assign n_19363 = ~n_19358 &  n_19362;
assign n_19364 =  n_18448 & ~n_19363;
assign n_19365 = ~n_19361 &  n_19364;
assign n_19366 = ~n_19353 & ~n_19365;
assign n_19367 =  n_19341 &  n_19366;
assign n_19368 =  x_503 & ~n_19367;
assign n_19369 = ~x_503 &  n_19367;
assign n_19370 = ~n_19368 & ~n_19369;
assign n_19371 = ~x_374 &  n_19323;
assign n_19372 =  x_374 & ~n_19323;
assign n_19373 = ~n_19371 & ~n_19372;
assign n_19374 = ~n_19327 & ~n_19331;
assign n_19375 =  n_19373 & ~n_19374;
assign n_19376 = ~n_19373 &  n_19374;
assign n_19377 = ~n_19375 & ~n_19376;
assign n_19378 = ~x_310 & ~n_19377;
assign n_19379 =  x_310 & ~n_19376;
assign n_19380 = ~n_19375 &  n_19379;
assign n_19381 =  n_18440 & ~n_19380;
assign n_19382 = ~n_19378 &  n_19381;
assign n_19383 =  x_502 & ~n_18431;
assign n_19384 =  x_1046 & ~n_19337;
assign n_19385 = ~x_1046 &  n_19337;
assign n_19386 =  n_18446 & ~n_19385;
assign n_19387 = ~n_19384 &  n_19386;
assign n_19388 = ~n_19383 & ~n_19387;
assign n_19389 = ~n_19382 &  n_19388;
assign n_19390 = ~x_118 &  n_19342;
assign n_19391 =  x_118 & ~n_19342;
assign n_19392 = ~n_19390 & ~n_19391;
assign n_19393 =  x_2839 & ~n_19348;
assign n_19394 = ~n_19347 & ~n_19393;
assign n_19395 =  n_19392 & ~n_19394;
assign n_19396 = ~n_19392 &  n_19394;
assign n_19397 = ~n_19395 & ~n_19396;
assign n_19398 = ~x_2838 & ~n_19397;
assign n_19399 =  x_2838 &  n_19397;
assign n_19400 =  n_18434 & ~n_19399;
assign n_19401 = ~n_19398 &  n_19400;
assign n_19402 = ~x_2038 &  n_19354;
assign n_19403 =  x_2038 & ~n_19354;
assign n_19404 = ~n_19402 & ~n_19403;
assign n_19405 = ~n_19358 & ~n_19362;
assign n_19406 =  n_19404 & ~n_19405;
assign n_19407 = ~n_19404 &  n_19405;
assign n_19408 = ~n_19406 & ~n_19407;
assign n_19409 = ~x_630 & ~n_19408;
assign n_19410 =  x_630 & ~n_19407;
assign n_19411 = ~n_19406 &  n_19410;
assign n_19412 =  n_18448 & ~n_19411;
assign n_19413 = ~n_19409 &  n_19412;
assign n_19414 = ~n_19401 & ~n_19413;
assign n_19415 =  n_19389 &  n_19414;
assign n_19416 =  x_502 & ~n_19415;
assign n_19417 = ~x_502 &  n_19415;
assign n_19418 = ~n_19416 & ~n_19417;
assign n_19419 = ~x_373 &  n_19371;
assign n_19420 =  x_373 & ~n_19371;
assign n_19421 = ~n_19419 & ~n_19420;
assign n_19422 = ~n_19375 & ~n_19379;
assign n_19423 =  n_19421 & ~n_19422;
assign n_19424 = ~n_19421 &  n_19422;
assign n_19425 = ~n_19423 & ~n_19424;
assign n_19426 = ~x_309 & ~n_19425;
assign n_19427 =  x_309 & ~n_19424;
assign n_19428 = ~n_19423 &  n_19427;
assign n_19429 =  n_18440 & ~n_19428;
assign n_19430 = ~n_19426 &  n_19429;
assign n_19431 =  x_501 & ~n_18431;
assign n_19432 =  x_1045 & ~n_19385;
assign n_19433 = ~x_1045 &  n_19385;
assign n_19434 =  n_18446 & ~n_19433;
assign n_19435 = ~n_19432 &  n_19434;
assign n_19436 = ~n_19431 & ~n_19435;
assign n_19437 = ~n_19430 &  n_19436;
assign n_19438 = ~x_117 &  n_19390;
assign n_19439 =  x_117 & ~n_19390;
assign n_19440 = ~n_19438 & ~n_19439;
assign n_19441 =  x_2838 & ~n_19396;
assign n_19442 = ~n_19395 & ~n_19441;
assign n_19443 =  n_19440 & ~n_19442;
assign n_19444 = ~n_19440 &  n_19442;
assign n_19445 = ~n_19443 & ~n_19444;
assign n_19446 = ~x_2837 & ~n_19445;
assign n_19447 =  x_2837 &  n_19445;
assign n_19448 =  n_18434 & ~n_19447;
assign n_19449 = ~n_19446 &  n_19448;
assign n_19450 = ~x_2037 &  n_19402;
assign n_19451 =  x_2037 & ~n_19402;
assign n_19452 = ~n_19450 & ~n_19451;
assign n_19453 = ~n_19406 & ~n_19410;
assign n_19454 =  n_19452 & ~n_19453;
assign n_19455 = ~n_19452 &  n_19453;
assign n_19456 = ~n_19454 & ~n_19455;
assign n_19457 = ~x_629 & ~n_19456;
assign n_19458 =  x_629 & ~n_19455;
assign n_19459 = ~n_19454 &  n_19458;
assign n_19460 =  n_18448 & ~n_19459;
assign n_19461 = ~n_19457 &  n_19460;
assign n_19462 = ~n_19449 & ~n_19461;
assign n_19463 =  n_19437 &  n_19462;
assign n_19464 =  x_501 & ~n_19463;
assign n_19465 = ~x_501 &  n_19463;
assign n_19466 = ~n_19464 & ~n_19465;
assign n_19467 = ~x_372 &  n_19419;
assign n_19468 =  x_372 & ~n_19419;
assign n_19469 = ~n_19467 & ~n_19468;
assign n_19470 = ~n_19423 & ~n_19427;
assign n_19471 =  n_19469 & ~n_19470;
assign n_19472 = ~n_19469 &  n_19470;
assign n_19473 = ~n_19471 & ~n_19472;
assign n_19474 = ~x_308 & ~n_19473;
assign n_19475 =  x_308 & ~n_19472;
assign n_19476 = ~n_19471 &  n_19475;
assign n_19477 =  n_18440 & ~n_19476;
assign n_19478 = ~n_19474 &  n_19477;
assign n_19479 =  x_500 & ~n_18431;
assign n_19480 =  x_1044 & ~n_19433;
assign n_19481 = ~x_1044 &  n_19433;
assign n_19482 =  n_18446 & ~n_19481;
assign n_19483 = ~n_19480 &  n_19482;
assign n_19484 = ~n_19479 & ~n_19483;
assign n_19485 = ~n_19478 &  n_19484;
assign n_19486 = ~x_116 &  n_19438;
assign n_19487 =  x_116 & ~n_19438;
assign n_19488 = ~n_19486 & ~n_19487;
assign n_19489 =  x_2837 & ~n_19444;
assign n_19490 = ~n_19443 & ~n_19489;
assign n_19491 =  n_19488 & ~n_19490;
assign n_19492 = ~n_19488 &  n_19490;
assign n_19493 = ~n_19491 & ~n_19492;
assign n_19494 = ~x_2836 & ~n_19493;
assign n_19495 =  x_2836 &  n_19493;
assign n_19496 =  n_18434 & ~n_19495;
assign n_19497 = ~n_19494 &  n_19496;
assign n_19498 = ~x_2036 &  n_19450;
assign n_19499 =  x_2036 & ~n_19450;
assign n_19500 = ~n_19498 & ~n_19499;
assign n_19501 = ~n_19454 & ~n_19458;
assign n_19502 =  n_19500 & ~n_19501;
assign n_19503 = ~n_19500 &  n_19501;
assign n_19504 = ~n_19502 & ~n_19503;
assign n_19505 = ~x_628 & ~n_19504;
assign n_19506 =  x_628 & ~n_19503;
assign n_19507 = ~n_19502 &  n_19506;
assign n_19508 =  n_18448 & ~n_19507;
assign n_19509 = ~n_19505 &  n_19508;
assign n_19510 = ~n_19497 & ~n_19509;
assign n_19511 =  n_19485 &  n_19510;
assign n_19512 =  x_500 & ~n_19511;
assign n_19513 = ~x_500 &  n_19511;
assign n_19514 = ~n_19512 & ~n_19513;
assign n_19515 = ~x_371 &  n_19467;
assign n_19516 =  x_371 & ~n_19467;
assign n_19517 = ~n_19515 & ~n_19516;
assign n_19518 = ~n_19471 & ~n_19475;
assign n_19519 =  n_19517 & ~n_19518;
assign n_19520 = ~n_19517 &  n_19518;
assign n_19521 = ~n_19519 & ~n_19520;
assign n_19522 = ~x_307 & ~n_19521;
assign n_19523 =  x_307 & ~n_19520;
assign n_19524 = ~n_19519 &  n_19523;
assign n_19525 =  n_18440 & ~n_19524;
assign n_19526 = ~n_19522 &  n_19525;
assign n_19527 =  x_499 & ~n_18431;
assign n_19528 =  x_1043 & ~n_19481;
assign n_19529 = ~x_1043 &  n_19481;
assign n_19530 =  n_18446 & ~n_19529;
assign n_19531 = ~n_19528 &  n_19530;
assign n_19532 = ~n_19527 & ~n_19531;
assign n_19533 = ~n_19526 &  n_19532;
assign n_19534 = ~x_115 &  n_19486;
assign n_19535 =  x_115 & ~n_19486;
assign n_19536 = ~n_19534 & ~n_19535;
assign n_19537 =  x_2836 & ~n_19492;
assign n_19538 = ~n_19491 & ~n_19537;
assign n_19539 =  n_19536 & ~n_19538;
assign n_19540 = ~n_19536 &  n_19538;
assign n_19541 = ~n_19539 & ~n_19540;
assign n_19542 = ~x_2835 & ~n_19541;
assign n_19543 =  x_2835 &  n_19541;
assign n_19544 =  n_18434 & ~n_19543;
assign n_19545 = ~n_19542 &  n_19544;
assign n_19546 = ~x_2035 &  n_19498;
assign n_19547 =  x_2035 & ~n_19498;
assign n_19548 = ~n_19546 & ~n_19547;
assign n_19549 = ~n_19502 & ~n_19506;
assign n_19550 =  n_19548 & ~n_19549;
assign n_19551 = ~n_19548 &  n_19549;
assign n_19552 = ~n_19550 & ~n_19551;
assign n_19553 = ~x_627 & ~n_19552;
assign n_19554 =  x_627 & ~n_19551;
assign n_19555 = ~n_19550 &  n_19554;
assign n_19556 =  n_18448 & ~n_19555;
assign n_19557 = ~n_19553 &  n_19556;
assign n_19558 = ~n_19545 & ~n_19557;
assign n_19559 =  n_19533 &  n_19558;
assign n_19560 =  x_499 & ~n_19559;
assign n_19561 = ~x_499 &  n_19559;
assign n_19562 = ~n_19560 & ~n_19561;
assign n_19563 = ~x_370 &  n_19515;
assign n_19564 =  x_370 & ~n_19515;
assign n_19565 = ~n_19563 & ~n_19564;
assign n_19566 = ~n_19519 & ~n_19523;
assign n_19567 =  n_19565 & ~n_19566;
assign n_19568 = ~n_19565 &  n_19566;
assign n_19569 = ~n_19567 & ~n_19568;
assign n_19570 = ~x_306 & ~n_19569;
assign n_19571 =  x_306 & ~n_19568;
assign n_19572 = ~n_19567 &  n_19571;
assign n_19573 =  n_18440 & ~n_19572;
assign n_19574 = ~n_19570 &  n_19573;
assign n_19575 =  x_498 & ~n_18431;
assign n_19576 =  x_1042 & ~n_19529;
assign n_19577 = ~x_1042 &  n_19529;
assign n_19578 =  n_18446 & ~n_19577;
assign n_19579 = ~n_19576 &  n_19578;
assign n_19580 = ~n_19575 & ~n_19579;
assign n_19581 = ~n_19574 &  n_19580;
assign n_19582 = ~x_114 &  n_19534;
assign n_19583 =  x_114 & ~n_19534;
assign n_19584 = ~n_19582 & ~n_19583;
assign n_19585 =  x_2835 & ~n_19540;
assign n_19586 = ~n_19539 & ~n_19585;
assign n_19587 =  n_19584 & ~n_19586;
assign n_19588 = ~n_19584 &  n_19586;
assign n_19589 = ~n_19587 & ~n_19588;
assign n_19590 = ~x_2834 & ~n_19589;
assign n_19591 =  x_2834 &  n_19589;
assign n_19592 =  n_18434 & ~n_19591;
assign n_19593 = ~n_19590 &  n_19592;
assign n_19594 = ~x_2034 &  n_19546;
assign n_19595 =  x_2034 & ~n_19546;
assign n_19596 = ~n_19594 & ~n_19595;
assign n_19597 = ~n_19550 & ~n_19554;
assign n_19598 =  n_19596 & ~n_19597;
assign n_19599 = ~n_19596 &  n_19597;
assign n_19600 = ~n_19598 & ~n_19599;
assign n_19601 = ~x_626 & ~n_19600;
assign n_19602 =  x_626 & ~n_19599;
assign n_19603 = ~n_19598 &  n_19602;
assign n_19604 =  n_18448 & ~n_19603;
assign n_19605 = ~n_19601 &  n_19604;
assign n_19606 = ~n_19593 & ~n_19605;
assign n_19607 =  n_19581 &  n_19606;
assign n_19608 =  x_498 & ~n_19607;
assign n_19609 = ~x_498 &  n_19607;
assign n_19610 = ~n_19608 & ~n_19609;
assign n_19611 = ~x_369 &  n_19563;
assign n_19612 =  x_369 & ~n_19563;
assign n_19613 = ~n_19611 & ~n_19612;
assign n_19614 = ~n_19567 & ~n_19571;
assign n_19615 =  n_19613 & ~n_19614;
assign n_19616 = ~n_19613 &  n_19614;
assign n_19617 = ~n_19615 & ~n_19616;
assign n_19618 = ~x_305 & ~n_19617;
assign n_19619 =  x_305 & ~n_19616;
assign n_19620 = ~n_19615 &  n_19619;
assign n_19621 =  n_18440 & ~n_19620;
assign n_19622 = ~n_19618 &  n_19621;
assign n_19623 =  x_497 & ~n_18431;
assign n_19624 =  x_1041 & ~n_19577;
assign n_19625 = ~x_1041 &  n_19577;
assign n_19626 =  n_18446 & ~n_19625;
assign n_19627 = ~n_19624 &  n_19626;
assign n_19628 = ~n_19623 & ~n_19627;
assign n_19629 = ~n_19622 &  n_19628;
assign n_19630 = ~x_113 &  n_19582;
assign n_19631 =  x_113 & ~n_19582;
assign n_19632 = ~n_19630 & ~n_19631;
assign n_19633 =  x_2834 & ~n_19588;
assign n_19634 = ~n_19587 & ~n_19633;
assign n_19635 =  n_19632 & ~n_19634;
assign n_19636 = ~n_19632 &  n_19634;
assign n_19637 = ~n_19635 & ~n_19636;
assign n_19638 = ~x_2833 & ~n_19637;
assign n_19639 =  x_2833 &  n_19637;
assign n_19640 =  n_18434 & ~n_19639;
assign n_19641 = ~n_19638 &  n_19640;
assign n_19642 = ~x_2033 &  n_19594;
assign n_19643 =  x_2033 & ~n_19594;
assign n_19644 = ~n_19642 & ~n_19643;
assign n_19645 = ~n_19598 & ~n_19602;
assign n_19646 =  n_19644 & ~n_19645;
assign n_19647 = ~n_19644 &  n_19645;
assign n_19648 = ~n_19646 & ~n_19647;
assign n_19649 = ~x_625 & ~n_19648;
assign n_19650 =  x_625 & ~n_19647;
assign n_19651 = ~n_19646 &  n_19650;
assign n_19652 =  n_18448 & ~n_19651;
assign n_19653 = ~n_19649 &  n_19652;
assign n_19654 = ~n_19641 & ~n_19653;
assign n_19655 =  n_19629 &  n_19654;
assign n_19656 =  x_497 & ~n_19655;
assign n_19657 = ~x_497 &  n_19655;
assign n_19658 = ~n_19656 & ~n_19657;
assign n_19659 = ~x_368 &  n_19611;
assign n_19660 =  x_368 & ~n_19611;
assign n_19661 = ~n_19659 & ~n_19660;
assign n_19662 = ~n_19615 & ~n_19619;
assign n_19663 =  n_19661 & ~n_19662;
assign n_19664 = ~n_19661 &  n_19662;
assign n_19665 = ~n_19663 & ~n_19664;
assign n_19666 = ~x_304 & ~n_19665;
assign n_19667 =  x_304 & ~n_19664;
assign n_19668 = ~n_19663 &  n_19667;
assign n_19669 =  n_18440 & ~n_19668;
assign n_19670 = ~n_19666 &  n_19669;
assign n_19671 =  x_496 & ~n_18431;
assign n_19672 =  x_1040 & ~n_19625;
assign n_19673 = ~x_1040 &  n_19625;
assign n_19674 =  n_18446 & ~n_19673;
assign n_19675 = ~n_19672 &  n_19674;
assign n_19676 = ~n_19671 & ~n_19675;
assign n_19677 = ~n_19670 &  n_19676;
assign n_19678 = ~x_112 &  n_19630;
assign n_19679 =  x_112 & ~n_19630;
assign n_19680 = ~n_19678 & ~n_19679;
assign n_19681 =  x_2833 & ~n_19636;
assign n_19682 = ~n_19635 & ~n_19681;
assign n_19683 =  n_19680 & ~n_19682;
assign n_19684 = ~n_19680 &  n_19682;
assign n_19685 = ~n_19683 & ~n_19684;
assign n_19686 = ~x_2832 & ~n_19685;
assign n_19687 =  x_2832 &  n_19685;
assign n_19688 =  n_18434 & ~n_19687;
assign n_19689 = ~n_19686 &  n_19688;
assign n_19690 = ~x_2032 &  n_19642;
assign n_19691 =  x_2032 & ~n_19642;
assign n_19692 = ~n_19690 & ~n_19691;
assign n_19693 = ~n_19646 & ~n_19650;
assign n_19694 =  n_19692 & ~n_19693;
assign n_19695 = ~n_19692 &  n_19693;
assign n_19696 = ~n_19694 & ~n_19695;
assign n_19697 = ~x_624 & ~n_19696;
assign n_19698 =  x_624 & ~n_19695;
assign n_19699 = ~n_19694 &  n_19698;
assign n_19700 =  n_18448 & ~n_19699;
assign n_19701 = ~n_19697 &  n_19700;
assign n_19702 = ~n_19689 & ~n_19701;
assign n_19703 =  n_19677 &  n_19702;
assign n_19704 =  x_496 & ~n_19703;
assign n_19705 = ~x_496 &  n_19703;
assign n_19706 = ~n_19704 & ~n_19705;
assign n_19707 = ~x_367 &  n_19659;
assign n_19708 =  x_367 & ~n_19659;
assign n_19709 = ~n_19707 & ~n_19708;
assign n_19710 = ~n_19663 & ~n_19667;
assign n_19711 =  n_19709 & ~n_19710;
assign n_19712 = ~n_19709 &  n_19710;
assign n_19713 = ~n_19711 & ~n_19712;
assign n_19714 = ~x_303 & ~n_19713;
assign n_19715 =  x_303 & ~n_19712;
assign n_19716 = ~n_19711 &  n_19715;
assign n_19717 =  n_18440 & ~n_19716;
assign n_19718 = ~n_19714 &  n_19717;
assign n_19719 =  x_495 & ~n_18431;
assign n_19720 =  x_1039 & ~n_19673;
assign n_19721 = ~x_1039 &  n_19673;
assign n_19722 =  n_18446 & ~n_19721;
assign n_19723 = ~n_19720 &  n_19722;
assign n_19724 = ~n_19719 & ~n_19723;
assign n_19725 = ~n_19718 &  n_19724;
assign n_19726 = ~x_111 &  n_19678;
assign n_19727 =  x_111 & ~n_19678;
assign n_19728 = ~n_19726 & ~n_19727;
assign n_19729 =  x_2832 & ~n_19684;
assign n_19730 = ~n_19683 & ~n_19729;
assign n_19731 =  n_19728 & ~n_19730;
assign n_19732 = ~n_19728 &  n_19730;
assign n_19733 = ~n_19731 & ~n_19732;
assign n_19734 = ~x_2831 & ~n_19733;
assign n_19735 =  x_2831 &  n_19733;
assign n_19736 =  n_18434 & ~n_19735;
assign n_19737 = ~n_19734 &  n_19736;
assign n_19738 = ~x_2031 &  n_19690;
assign n_19739 =  x_2031 & ~n_19690;
assign n_19740 = ~n_19738 & ~n_19739;
assign n_19741 = ~n_19694 & ~n_19698;
assign n_19742 =  n_19740 & ~n_19741;
assign n_19743 = ~n_19740 &  n_19741;
assign n_19744 = ~n_19742 & ~n_19743;
assign n_19745 = ~x_623 & ~n_19744;
assign n_19746 =  x_623 & ~n_19743;
assign n_19747 = ~n_19742 &  n_19746;
assign n_19748 =  n_18448 & ~n_19747;
assign n_19749 = ~n_19745 &  n_19748;
assign n_19750 = ~n_19737 & ~n_19749;
assign n_19751 =  n_19725 &  n_19750;
assign n_19752 =  x_495 & ~n_19751;
assign n_19753 = ~x_495 &  n_19751;
assign n_19754 = ~n_19752 & ~n_19753;
assign n_19755 = ~x_366 &  n_19707;
assign n_19756 =  x_366 & ~n_19707;
assign n_19757 = ~n_19755 & ~n_19756;
assign n_19758 = ~n_19711 & ~n_19715;
assign n_19759 =  n_19757 & ~n_19758;
assign n_19760 = ~n_19757 &  n_19758;
assign n_19761 = ~n_19759 & ~n_19760;
assign n_19762 = ~x_302 & ~n_19761;
assign n_19763 =  x_302 & ~n_19760;
assign n_19764 = ~n_19759 &  n_19763;
assign n_19765 =  n_18440 & ~n_19764;
assign n_19766 = ~n_19762 &  n_19765;
assign n_19767 =  x_494 & ~n_18431;
assign n_19768 =  x_1038 & ~n_19721;
assign n_19769 = ~x_1038 &  n_19721;
assign n_19770 =  n_18446 & ~n_19769;
assign n_19771 = ~n_19768 &  n_19770;
assign n_19772 = ~n_19767 & ~n_19771;
assign n_19773 = ~n_19766 &  n_19772;
assign n_19774 = ~x_110 &  n_19726;
assign n_19775 =  x_110 & ~n_19726;
assign n_19776 = ~n_19774 & ~n_19775;
assign n_19777 =  x_2831 & ~n_19732;
assign n_19778 = ~n_19731 & ~n_19777;
assign n_19779 =  n_19776 & ~n_19778;
assign n_19780 = ~n_19776 &  n_19778;
assign n_19781 = ~n_19779 & ~n_19780;
assign n_19782 = ~x_2830 & ~n_19781;
assign n_19783 =  x_2830 &  n_19781;
assign n_19784 =  n_18434 & ~n_19783;
assign n_19785 = ~n_19782 &  n_19784;
assign n_19786 = ~x_2030 &  n_19738;
assign n_19787 =  x_2030 & ~n_19738;
assign n_19788 = ~n_19786 & ~n_19787;
assign n_19789 = ~n_19742 & ~n_19746;
assign n_19790 =  n_19788 & ~n_19789;
assign n_19791 = ~n_19788 &  n_19789;
assign n_19792 = ~n_19790 & ~n_19791;
assign n_19793 = ~x_622 & ~n_19792;
assign n_19794 =  x_622 & ~n_19791;
assign n_19795 = ~n_19790 &  n_19794;
assign n_19796 =  n_18448 & ~n_19795;
assign n_19797 = ~n_19793 &  n_19796;
assign n_19798 = ~n_19785 & ~n_19797;
assign n_19799 =  n_19773 &  n_19798;
assign n_19800 =  x_494 & ~n_19799;
assign n_19801 = ~x_494 &  n_19799;
assign n_19802 = ~n_19800 & ~n_19801;
assign n_19803 = ~x_365 &  n_19755;
assign n_19804 =  x_365 & ~n_19755;
assign n_19805 = ~n_19803 & ~n_19804;
assign n_19806 = ~n_19759 & ~n_19763;
assign n_19807 =  n_19805 & ~n_19806;
assign n_19808 = ~n_19805 &  n_19806;
assign n_19809 = ~n_19807 & ~n_19808;
assign n_19810 = ~x_301 & ~n_19809;
assign n_19811 =  x_301 & ~n_19808;
assign n_19812 = ~n_19807 &  n_19811;
assign n_19813 =  n_18440 & ~n_19812;
assign n_19814 = ~n_19810 &  n_19813;
assign n_19815 =  x_493 & ~n_18431;
assign n_19816 =  x_1037 & ~n_19769;
assign n_19817 = ~x_1037 &  n_19769;
assign n_19818 =  n_18446 & ~n_19817;
assign n_19819 = ~n_19816 &  n_19818;
assign n_19820 = ~n_19815 & ~n_19819;
assign n_19821 = ~n_19814 &  n_19820;
assign n_19822 = ~x_109 &  n_19774;
assign n_19823 =  x_109 & ~n_19774;
assign n_19824 = ~n_19822 & ~n_19823;
assign n_19825 =  x_2830 & ~n_19780;
assign n_19826 = ~n_19779 & ~n_19825;
assign n_19827 =  n_19824 & ~n_19826;
assign n_19828 = ~n_19824 &  n_19826;
assign n_19829 = ~n_19827 & ~n_19828;
assign n_19830 = ~x_2829 & ~n_19829;
assign n_19831 =  x_2829 &  n_19829;
assign n_19832 =  n_18434 & ~n_19831;
assign n_19833 = ~n_19830 &  n_19832;
assign n_19834 = ~x_2029 &  n_19786;
assign n_19835 =  x_2029 & ~n_19786;
assign n_19836 = ~n_19834 & ~n_19835;
assign n_19837 = ~n_19790 & ~n_19794;
assign n_19838 =  n_19836 & ~n_19837;
assign n_19839 = ~n_19836 &  n_19837;
assign n_19840 = ~n_19838 & ~n_19839;
assign n_19841 = ~x_621 & ~n_19840;
assign n_19842 =  x_621 & ~n_19839;
assign n_19843 = ~n_19838 &  n_19842;
assign n_19844 =  n_18448 & ~n_19843;
assign n_19845 = ~n_19841 &  n_19844;
assign n_19846 = ~n_19833 & ~n_19845;
assign n_19847 =  n_19821 &  n_19846;
assign n_19848 =  x_493 & ~n_19847;
assign n_19849 = ~x_493 &  n_19847;
assign n_19850 = ~n_19848 & ~n_19849;
assign n_19851 = ~x_364 &  n_19803;
assign n_19852 =  x_364 & ~n_19803;
assign n_19853 = ~n_19851 & ~n_19852;
assign n_19854 = ~n_19807 & ~n_19811;
assign n_19855 =  n_19853 & ~n_19854;
assign n_19856 = ~n_19853 &  n_19854;
assign n_19857 = ~n_19855 & ~n_19856;
assign n_19858 = ~x_300 & ~n_19857;
assign n_19859 =  x_300 & ~n_19856;
assign n_19860 = ~n_19855 &  n_19859;
assign n_19861 =  n_18440 & ~n_19860;
assign n_19862 = ~n_19858 &  n_19861;
assign n_19863 =  x_492 & ~n_18431;
assign n_19864 =  x_1036 & ~n_19817;
assign n_19865 = ~x_1036 &  n_19817;
assign n_19866 =  n_18446 & ~n_19865;
assign n_19867 = ~n_19864 &  n_19866;
assign n_19868 = ~n_19863 & ~n_19867;
assign n_19869 = ~n_19862 &  n_19868;
assign n_19870 = ~x_108 &  n_19822;
assign n_19871 =  x_108 & ~n_19822;
assign n_19872 = ~n_19870 & ~n_19871;
assign n_19873 =  x_2829 & ~n_19828;
assign n_19874 = ~n_19827 & ~n_19873;
assign n_19875 =  n_19872 & ~n_19874;
assign n_19876 = ~n_19872 &  n_19874;
assign n_19877 = ~n_19875 & ~n_19876;
assign n_19878 = ~x_2828 & ~n_19877;
assign n_19879 =  x_2828 &  n_19877;
assign n_19880 =  n_18434 & ~n_19879;
assign n_19881 = ~n_19878 &  n_19880;
assign n_19882 = ~x_2028 &  n_19834;
assign n_19883 =  x_2028 & ~n_19834;
assign n_19884 = ~n_19882 & ~n_19883;
assign n_19885 = ~n_19838 & ~n_19842;
assign n_19886 =  n_19884 & ~n_19885;
assign n_19887 = ~n_19884 &  n_19885;
assign n_19888 = ~n_19886 & ~n_19887;
assign n_19889 = ~x_620 & ~n_19888;
assign n_19890 =  x_620 & ~n_19887;
assign n_19891 = ~n_19886 &  n_19890;
assign n_19892 =  n_18448 & ~n_19891;
assign n_19893 = ~n_19889 &  n_19892;
assign n_19894 = ~n_19881 & ~n_19893;
assign n_19895 =  n_19869 &  n_19894;
assign n_19896 =  x_492 & ~n_19895;
assign n_19897 = ~x_492 &  n_19895;
assign n_19898 = ~n_19896 & ~n_19897;
assign n_19899 =  x_2828 & ~n_19876;
assign n_19900 = ~n_19875 & ~n_19899;
assign n_19901 =  x_107 & ~x_2827;
assign n_19902 = ~x_107 &  x_2827;
assign n_19903 = ~n_19901 & ~n_19902;
assign n_19904 =  n_19870 &  n_19903;
assign n_19905 = ~n_19870 & ~n_19903;
assign n_19906 = ~n_19904 & ~n_19905;
assign n_19907 = ~n_19900 &  n_19906;
assign n_19908 =  n_19900 & ~n_19906;
assign n_19909 =  n_18434 & ~n_19908;
assign n_19910 = ~n_19907 &  n_19909;
assign n_19911 =  x_491 & ~n_18431;
assign n_19912 = ~x_1035 &  n_19865;
assign n_19913 =  x_1035 & ~n_19865;
assign n_19914 =  n_18446 & ~n_19913;
assign n_19915 = ~n_19912 &  n_19914;
assign n_19916 = ~n_19911 & ~n_19915;
assign n_19917 = ~n_19910 &  n_19916;
assign n_19918 = ~n_19886 & ~n_19890;
assign n_19919 =  x_619 & ~x_2027;
assign n_19920 = ~x_619 &  x_2027;
assign n_19921 = ~n_19919 & ~n_19920;
assign n_19922 =  n_19882 &  n_19921;
assign n_19923 = ~n_19882 & ~n_19921;
assign n_19924 = ~n_19922 & ~n_19923;
assign n_19925 =  n_19918 & ~n_19924;
assign n_19926 = ~n_19918 &  n_19924;
assign n_19927 =  n_18448 & ~n_19926;
assign n_19928 = ~n_19925 &  n_19927;
assign n_19929 = ~n_19855 & ~n_19859;
assign n_19930 =  x_299 & ~x_363;
assign n_19931 = ~x_299 &  x_363;
assign n_19932 = ~n_19930 & ~n_19931;
assign n_19933 =  n_19851 &  n_19932;
assign n_19934 = ~n_19851 & ~n_19932;
assign n_19935 = ~n_19933 & ~n_19934;
assign n_19936 =  n_19929 & ~n_19935;
assign n_19937 = ~n_19929 &  n_19935;
assign n_19938 =  n_18440 & ~n_19937;
assign n_19939 = ~n_19936 &  n_19938;
assign n_19940 = ~n_19928 & ~n_19939;
assign n_19941 =  n_19917 &  n_19940;
assign n_19942 =  x_491 & ~n_19941;
assign n_19943 = ~x_491 &  n_19941;
assign n_19944 = ~n_19942 & ~n_19943;
assign n_19945 =  n_2 &  n_2886;
assign n_19946 =  n_19945 &  n_3860;
assign n_19947 =  x_490 & ~n_19946;
assign n_19948 =  i_32 &  n_19946;
assign n_19949 = ~n_19947 & ~n_19948;
assign n_19950 =  x_490 & ~n_19949;
assign n_19951 = ~x_490 &  n_19949;
assign n_19952 = ~n_19950 & ~n_19951;
assign n_19953 =  x_489 & ~n_19946;
assign n_19954 =  i_31 &  n_19946;
assign n_19955 = ~n_19953 & ~n_19954;
assign n_19956 =  x_489 & ~n_19955;
assign n_19957 = ~x_489 &  n_19955;
assign n_19958 = ~n_19956 & ~n_19957;
assign n_19959 =  x_488 & ~n_19946;
assign n_19960 =  i_30 &  n_19946;
assign n_19961 = ~n_19959 & ~n_19960;
assign n_19962 =  x_488 & ~n_19961;
assign n_19963 = ~x_488 &  n_19961;
assign n_19964 = ~n_19962 & ~n_19963;
assign n_19965 =  x_487 & ~n_19946;
assign n_19966 =  i_29 &  n_19946;
assign n_19967 = ~n_19965 & ~n_19966;
assign n_19968 =  x_487 & ~n_19967;
assign n_19969 = ~x_487 &  n_19967;
assign n_19970 = ~n_19968 & ~n_19969;
assign n_19971 =  x_486 & ~n_19946;
assign n_19972 =  i_28 &  n_19946;
assign n_19973 = ~n_19971 & ~n_19972;
assign n_19974 =  x_486 & ~n_19973;
assign n_19975 = ~x_486 &  n_19973;
assign n_19976 = ~n_19974 & ~n_19975;
assign n_19977 =  x_485 & ~n_19946;
assign n_19978 =  i_27 &  n_19946;
assign n_19979 = ~n_19977 & ~n_19978;
assign n_19980 =  x_485 & ~n_19979;
assign n_19981 = ~x_485 &  n_19979;
assign n_19982 = ~n_19980 & ~n_19981;
assign n_19983 =  x_484 & ~n_19946;
assign n_19984 =  i_26 &  n_19946;
assign n_19985 = ~n_19983 & ~n_19984;
assign n_19986 =  x_484 & ~n_19985;
assign n_19987 = ~x_484 &  n_19985;
assign n_19988 = ~n_19986 & ~n_19987;
assign n_19989 =  x_483 & ~n_19946;
assign n_19990 =  i_25 &  n_19946;
assign n_19991 = ~n_19989 & ~n_19990;
assign n_19992 =  x_483 & ~n_19991;
assign n_19993 = ~x_483 &  n_19991;
assign n_19994 = ~n_19992 & ~n_19993;
assign n_19995 =  x_482 & ~n_19946;
assign n_19996 =  i_24 &  n_19946;
assign n_19997 = ~n_19995 & ~n_19996;
assign n_19998 =  x_482 & ~n_19997;
assign n_19999 = ~x_482 &  n_19997;
assign n_20000 = ~n_19998 & ~n_19999;
assign n_20001 =  x_481 & ~n_19946;
assign n_20002 =  i_23 &  n_19946;
assign n_20003 = ~n_20001 & ~n_20002;
assign n_20004 =  x_481 & ~n_20003;
assign n_20005 = ~x_481 &  n_20003;
assign n_20006 = ~n_20004 & ~n_20005;
assign n_20007 =  x_480 & ~n_19946;
assign n_20008 =  i_22 &  n_19946;
assign n_20009 = ~n_20007 & ~n_20008;
assign n_20010 =  x_480 & ~n_20009;
assign n_20011 = ~x_480 &  n_20009;
assign n_20012 = ~n_20010 & ~n_20011;
assign n_20013 =  x_479 & ~n_19946;
assign n_20014 =  i_21 &  n_19946;
assign n_20015 = ~n_20013 & ~n_20014;
assign n_20016 =  x_479 & ~n_20015;
assign n_20017 = ~x_479 &  n_20015;
assign n_20018 = ~n_20016 & ~n_20017;
assign n_20019 =  x_478 & ~n_19946;
assign n_20020 =  i_20 &  n_19946;
assign n_20021 = ~n_20019 & ~n_20020;
assign n_20022 =  x_478 & ~n_20021;
assign n_20023 = ~x_478 &  n_20021;
assign n_20024 = ~n_20022 & ~n_20023;
assign n_20025 =  x_477 & ~n_19946;
assign n_20026 =  i_19 &  n_19946;
assign n_20027 = ~n_20025 & ~n_20026;
assign n_20028 =  x_477 & ~n_20027;
assign n_20029 = ~x_477 &  n_20027;
assign n_20030 = ~n_20028 & ~n_20029;
assign n_20031 =  x_476 & ~n_19946;
assign n_20032 =  i_18 &  n_19946;
assign n_20033 = ~n_20031 & ~n_20032;
assign n_20034 =  x_476 & ~n_20033;
assign n_20035 = ~x_476 &  n_20033;
assign n_20036 = ~n_20034 & ~n_20035;
assign n_20037 =  x_475 & ~n_19946;
assign n_20038 =  i_17 &  n_19946;
assign n_20039 = ~n_20037 & ~n_20038;
assign n_20040 =  x_475 & ~n_20039;
assign n_20041 = ~x_475 &  n_20039;
assign n_20042 = ~n_20040 & ~n_20041;
assign n_20043 =  x_474 & ~n_19946;
assign n_20044 =  i_16 &  n_19946;
assign n_20045 = ~n_20043 & ~n_20044;
assign n_20046 =  x_474 & ~n_20045;
assign n_20047 = ~x_474 &  n_20045;
assign n_20048 = ~n_20046 & ~n_20047;
assign n_20049 =  x_473 & ~n_19946;
assign n_20050 =  i_15 &  n_19946;
assign n_20051 = ~n_20049 & ~n_20050;
assign n_20052 =  x_473 & ~n_20051;
assign n_20053 = ~x_473 &  n_20051;
assign n_20054 = ~n_20052 & ~n_20053;
assign n_20055 =  x_472 & ~n_19946;
assign n_20056 =  i_14 &  n_19946;
assign n_20057 = ~n_20055 & ~n_20056;
assign n_20058 =  x_472 & ~n_20057;
assign n_20059 = ~x_472 &  n_20057;
assign n_20060 = ~n_20058 & ~n_20059;
assign n_20061 =  x_471 & ~n_19946;
assign n_20062 =  i_13 &  n_19946;
assign n_20063 = ~n_20061 & ~n_20062;
assign n_20064 =  x_471 & ~n_20063;
assign n_20065 = ~x_471 &  n_20063;
assign n_20066 = ~n_20064 & ~n_20065;
assign n_20067 =  x_470 & ~n_19946;
assign n_20068 =  i_12 &  n_19946;
assign n_20069 = ~n_20067 & ~n_20068;
assign n_20070 =  x_470 & ~n_20069;
assign n_20071 = ~x_470 &  n_20069;
assign n_20072 = ~n_20070 & ~n_20071;
assign n_20073 =  x_469 & ~n_19946;
assign n_20074 =  i_11 &  n_19946;
assign n_20075 = ~n_20073 & ~n_20074;
assign n_20076 =  x_469 & ~n_20075;
assign n_20077 = ~x_469 &  n_20075;
assign n_20078 = ~n_20076 & ~n_20077;
assign n_20079 =  x_468 & ~n_19946;
assign n_20080 =  i_10 &  n_19946;
assign n_20081 = ~n_20079 & ~n_20080;
assign n_20082 =  x_468 & ~n_20081;
assign n_20083 = ~x_468 &  n_20081;
assign n_20084 = ~n_20082 & ~n_20083;
assign n_20085 =  x_467 & ~n_19946;
assign n_20086 =  i_9 &  n_19946;
assign n_20087 = ~n_20085 & ~n_20086;
assign n_20088 =  x_467 & ~n_20087;
assign n_20089 = ~x_467 &  n_20087;
assign n_20090 = ~n_20088 & ~n_20089;
assign n_20091 =  x_466 & ~n_19946;
assign n_20092 =  i_8 &  n_19946;
assign n_20093 = ~n_20091 & ~n_20092;
assign n_20094 =  x_466 & ~n_20093;
assign n_20095 = ~x_466 &  n_20093;
assign n_20096 = ~n_20094 & ~n_20095;
assign n_20097 =  x_465 & ~n_19946;
assign n_20098 =  i_7 &  n_19946;
assign n_20099 = ~n_20097 & ~n_20098;
assign n_20100 =  x_465 & ~n_20099;
assign n_20101 = ~x_465 &  n_20099;
assign n_20102 = ~n_20100 & ~n_20101;
assign n_20103 =  x_464 & ~n_19946;
assign n_20104 =  i_6 &  n_19946;
assign n_20105 = ~n_20103 & ~n_20104;
assign n_20106 =  x_464 & ~n_20105;
assign n_20107 = ~x_464 &  n_20105;
assign n_20108 = ~n_20106 & ~n_20107;
assign n_20109 =  x_463 & ~n_19946;
assign n_20110 =  i_5 &  n_19946;
assign n_20111 = ~n_20109 & ~n_20110;
assign n_20112 =  x_463 & ~n_20111;
assign n_20113 = ~x_463 &  n_20111;
assign n_20114 = ~n_20112 & ~n_20113;
assign n_20115 =  x_462 & ~n_19946;
assign n_20116 =  i_4 &  n_19946;
assign n_20117 = ~n_20115 & ~n_20116;
assign n_20118 =  x_462 & ~n_20117;
assign n_20119 = ~x_462 &  n_20117;
assign n_20120 = ~n_20118 & ~n_20119;
assign n_20121 =  x_461 & ~n_19946;
assign n_20122 =  i_3 &  n_19946;
assign n_20123 = ~n_20121 & ~n_20122;
assign n_20124 =  x_461 & ~n_20123;
assign n_20125 = ~x_461 &  n_20123;
assign n_20126 = ~n_20124 & ~n_20125;
assign n_20127 =  x_460 & ~n_19946;
assign n_20128 =  i_2 &  n_19946;
assign n_20129 = ~n_20127 & ~n_20128;
assign n_20130 =  x_460 & ~n_20129;
assign n_20131 = ~x_460 &  n_20129;
assign n_20132 = ~n_20130 & ~n_20131;
assign n_20133 =  x_459 & ~n_19946;
assign n_20134 =  i_1 &  n_19946;
assign n_20135 = ~n_20133 & ~n_20134;
assign n_20136 =  x_459 & ~n_20135;
assign n_20137 = ~x_459 &  n_20135;
assign n_20138 = ~n_20136 & ~n_20137;
assign n_20139 =  n_4993 &  n_191;
assign n_20140 =  x_458 & ~n_20139;
assign n_20141 =  i_32 &  n_20139;
assign n_20142 = ~n_20140 & ~n_20141;
assign n_20143 =  x_458 & ~n_20142;
assign n_20144 = ~x_458 &  n_20142;
assign n_20145 = ~n_20143 & ~n_20144;
assign n_20146 =  x_457 & ~n_20139;
assign n_20147 =  i_31 &  n_20139;
assign n_20148 = ~n_20146 & ~n_20147;
assign n_20149 =  x_457 & ~n_20148;
assign n_20150 = ~x_457 &  n_20148;
assign n_20151 = ~n_20149 & ~n_20150;
assign n_20152 =  x_456 & ~n_20139;
assign n_20153 =  i_30 &  n_20139;
assign n_20154 = ~n_20152 & ~n_20153;
assign n_20155 =  x_456 & ~n_20154;
assign n_20156 = ~x_456 &  n_20154;
assign n_20157 = ~n_20155 & ~n_20156;
assign n_20158 =  x_455 & ~n_20139;
assign n_20159 =  i_29 &  n_20139;
assign n_20160 = ~n_20158 & ~n_20159;
assign n_20161 =  x_455 & ~n_20160;
assign n_20162 = ~x_455 &  n_20160;
assign n_20163 = ~n_20161 & ~n_20162;
assign n_20164 =  x_454 & ~n_20139;
assign n_20165 =  i_28 &  n_20139;
assign n_20166 = ~n_20164 & ~n_20165;
assign n_20167 =  x_454 & ~n_20166;
assign n_20168 = ~x_454 &  n_20166;
assign n_20169 = ~n_20167 & ~n_20168;
assign n_20170 =  x_453 & ~n_20139;
assign n_20171 =  i_27 &  n_20139;
assign n_20172 = ~n_20170 & ~n_20171;
assign n_20173 =  x_453 & ~n_20172;
assign n_20174 = ~x_453 &  n_20172;
assign n_20175 = ~n_20173 & ~n_20174;
assign n_20176 =  x_452 & ~n_20139;
assign n_20177 =  i_26 &  n_20139;
assign n_20178 = ~n_20176 & ~n_20177;
assign n_20179 =  x_452 & ~n_20178;
assign n_20180 = ~x_452 &  n_20178;
assign n_20181 = ~n_20179 & ~n_20180;
assign n_20182 =  x_451 & ~n_20139;
assign n_20183 =  i_25 &  n_20139;
assign n_20184 = ~n_20182 & ~n_20183;
assign n_20185 =  x_451 & ~n_20184;
assign n_20186 = ~x_451 &  n_20184;
assign n_20187 = ~n_20185 & ~n_20186;
assign n_20188 =  x_450 & ~n_20139;
assign n_20189 =  i_24 &  n_20139;
assign n_20190 = ~n_20188 & ~n_20189;
assign n_20191 =  x_450 & ~n_20190;
assign n_20192 = ~x_450 &  n_20190;
assign n_20193 = ~n_20191 & ~n_20192;
assign n_20194 =  x_449 & ~n_20139;
assign n_20195 =  i_23 &  n_20139;
assign n_20196 = ~n_20194 & ~n_20195;
assign n_20197 =  x_449 & ~n_20196;
assign n_20198 = ~x_449 &  n_20196;
assign n_20199 = ~n_20197 & ~n_20198;
assign n_20200 =  x_448 & ~n_20139;
assign n_20201 =  i_22 &  n_20139;
assign n_20202 = ~n_20200 & ~n_20201;
assign n_20203 =  x_448 & ~n_20202;
assign n_20204 = ~x_448 &  n_20202;
assign n_20205 = ~n_20203 & ~n_20204;
assign n_20206 =  x_447 & ~n_20139;
assign n_20207 =  i_21 &  n_20139;
assign n_20208 = ~n_20206 & ~n_20207;
assign n_20209 =  x_447 & ~n_20208;
assign n_20210 = ~x_447 &  n_20208;
assign n_20211 = ~n_20209 & ~n_20210;
assign n_20212 =  x_446 & ~n_20139;
assign n_20213 =  i_20 &  n_20139;
assign n_20214 = ~n_20212 & ~n_20213;
assign n_20215 =  x_446 & ~n_20214;
assign n_20216 = ~x_446 &  n_20214;
assign n_20217 = ~n_20215 & ~n_20216;
assign n_20218 =  x_445 & ~n_20139;
assign n_20219 =  i_19 &  n_20139;
assign n_20220 = ~n_20218 & ~n_20219;
assign n_20221 =  x_445 & ~n_20220;
assign n_20222 = ~x_445 &  n_20220;
assign n_20223 = ~n_20221 & ~n_20222;
assign n_20224 =  x_444 & ~n_20139;
assign n_20225 =  i_18 &  n_20139;
assign n_20226 = ~n_20224 & ~n_20225;
assign n_20227 =  x_444 & ~n_20226;
assign n_20228 = ~x_444 &  n_20226;
assign n_20229 = ~n_20227 & ~n_20228;
assign n_20230 =  x_443 & ~n_20139;
assign n_20231 =  i_17 &  n_20139;
assign n_20232 = ~n_20230 & ~n_20231;
assign n_20233 =  x_443 & ~n_20232;
assign n_20234 = ~x_443 &  n_20232;
assign n_20235 = ~n_20233 & ~n_20234;
assign n_20236 =  x_442 & ~n_20139;
assign n_20237 =  i_16 &  n_20139;
assign n_20238 = ~n_20236 & ~n_20237;
assign n_20239 =  x_442 & ~n_20238;
assign n_20240 = ~x_442 &  n_20238;
assign n_20241 = ~n_20239 & ~n_20240;
assign n_20242 =  x_441 & ~n_20139;
assign n_20243 =  i_15 &  n_20139;
assign n_20244 = ~n_20242 & ~n_20243;
assign n_20245 =  x_441 & ~n_20244;
assign n_20246 = ~x_441 &  n_20244;
assign n_20247 = ~n_20245 & ~n_20246;
assign n_20248 =  x_440 & ~n_20139;
assign n_20249 =  i_14 &  n_20139;
assign n_20250 = ~n_20248 & ~n_20249;
assign n_20251 =  x_440 & ~n_20250;
assign n_20252 = ~x_440 &  n_20250;
assign n_20253 = ~n_20251 & ~n_20252;
assign n_20254 =  x_439 & ~n_20139;
assign n_20255 =  i_13 &  n_20139;
assign n_20256 = ~n_20254 & ~n_20255;
assign n_20257 =  x_439 & ~n_20256;
assign n_20258 = ~x_439 &  n_20256;
assign n_20259 = ~n_20257 & ~n_20258;
assign n_20260 =  x_438 & ~n_20139;
assign n_20261 =  i_12 &  n_20139;
assign n_20262 = ~n_20260 & ~n_20261;
assign n_20263 =  x_438 & ~n_20262;
assign n_20264 = ~x_438 &  n_20262;
assign n_20265 = ~n_20263 & ~n_20264;
assign n_20266 =  x_437 & ~n_20139;
assign n_20267 =  i_11 &  n_20139;
assign n_20268 = ~n_20266 & ~n_20267;
assign n_20269 =  x_437 & ~n_20268;
assign n_20270 = ~x_437 &  n_20268;
assign n_20271 = ~n_20269 & ~n_20270;
assign n_20272 =  x_436 & ~n_20139;
assign n_20273 =  i_10 &  n_20139;
assign n_20274 = ~n_20272 & ~n_20273;
assign n_20275 =  x_436 & ~n_20274;
assign n_20276 = ~x_436 &  n_20274;
assign n_20277 = ~n_20275 & ~n_20276;
assign n_20278 =  x_435 & ~n_20139;
assign n_20279 =  i_9 &  n_20139;
assign n_20280 = ~n_20278 & ~n_20279;
assign n_20281 =  x_435 & ~n_20280;
assign n_20282 = ~x_435 &  n_20280;
assign n_20283 = ~n_20281 & ~n_20282;
assign n_20284 =  x_434 & ~n_20139;
assign n_20285 =  i_8 &  n_20139;
assign n_20286 = ~n_20284 & ~n_20285;
assign n_20287 =  x_434 & ~n_20286;
assign n_20288 = ~x_434 &  n_20286;
assign n_20289 = ~n_20287 & ~n_20288;
assign n_20290 =  x_433 & ~n_20139;
assign n_20291 =  i_7 &  n_20139;
assign n_20292 = ~n_20290 & ~n_20291;
assign n_20293 =  x_433 & ~n_20292;
assign n_20294 = ~x_433 &  n_20292;
assign n_20295 = ~n_20293 & ~n_20294;
assign n_20296 =  x_432 & ~n_20139;
assign n_20297 =  i_6 &  n_20139;
assign n_20298 = ~n_20296 & ~n_20297;
assign n_20299 =  x_432 & ~n_20298;
assign n_20300 = ~x_432 &  n_20298;
assign n_20301 = ~n_20299 & ~n_20300;
assign n_20302 =  x_431 & ~n_20139;
assign n_20303 =  i_5 &  n_20139;
assign n_20304 = ~n_20302 & ~n_20303;
assign n_20305 =  x_431 & ~n_20304;
assign n_20306 = ~x_431 &  n_20304;
assign n_20307 = ~n_20305 & ~n_20306;
assign n_20308 =  x_430 & ~n_20139;
assign n_20309 =  i_4 &  n_20139;
assign n_20310 = ~n_20308 & ~n_20309;
assign n_20311 =  x_430 & ~n_20310;
assign n_20312 = ~x_430 &  n_20310;
assign n_20313 = ~n_20311 & ~n_20312;
assign n_20314 =  x_429 & ~n_20139;
assign n_20315 =  i_3 &  n_20139;
assign n_20316 = ~n_20314 & ~n_20315;
assign n_20317 =  x_429 & ~n_20316;
assign n_20318 = ~x_429 &  n_20316;
assign n_20319 = ~n_20317 & ~n_20318;
assign n_20320 =  x_428 & ~n_20139;
assign n_20321 =  i_2 &  n_20139;
assign n_20322 = ~n_20320 & ~n_20321;
assign n_20323 =  x_428 & ~n_20322;
assign n_20324 = ~x_428 &  n_20322;
assign n_20325 = ~n_20323 & ~n_20324;
assign n_20326 =  x_427 & ~n_20139;
assign n_20327 =  i_1 &  n_20139;
assign n_20328 = ~n_20326 & ~n_20327;
assign n_20329 =  x_427 & ~n_20328;
assign n_20330 = ~x_427 &  n_20328;
assign n_20331 = ~n_20329 & ~n_20330;
assign n_20332 =  n_2 &  n_12032;
assign n_20333 =  x_426 & ~n_20332;
assign n_20334 =  x_106 &  n_20332;
assign n_20335 = ~n_20333 & ~n_20334;
assign n_20336 =  x_426 & ~n_20335;
assign n_20337 = ~x_426 &  n_20335;
assign n_20338 = ~n_20336 & ~n_20337;
assign n_20339 =  x_425 & ~n_20332;
assign n_20340 =  x_105 &  n_20332;
assign n_20341 = ~n_20339 & ~n_20340;
assign n_20342 =  x_425 & ~n_20341;
assign n_20343 = ~x_425 &  n_20341;
assign n_20344 = ~n_20342 & ~n_20343;
assign n_20345 =  x_424 & ~n_20332;
assign n_20346 =  x_104 &  n_20332;
assign n_20347 = ~n_20345 & ~n_20346;
assign n_20348 =  x_424 & ~n_20347;
assign n_20349 = ~x_424 &  n_20347;
assign n_20350 = ~n_20348 & ~n_20349;
assign n_20351 =  x_423 & ~n_20332;
assign n_20352 =  x_103 &  n_20332;
assign n_20353 = ~n_20351 & ~n_20352;
assign n_20354 =  x_423 & ~n_20353;
assign n_20355 = ~x_423 &  n_20353;
assign n_20356 = ~n_20354 & ~n_20355;
assign n_20357 =  x_422 & ~n_20332;
assign n_20358 =  x_102 &  n_20332;
assign n_20359 = ~n_20357 & ~n_20358;
assign n_20360 =  x_422 & ~n_20359;
assign n_20361 = ~x_422 &  n_20359;
assign n_20362 = ~n_20360 & ~n_20361;
assign n_20363 =  x_421 & ~n_20332;
assign n_20364 =  x_101 &  n_20332;
assign n_20365 = ~n_20363 & ~n_20364;
assign n_20366 =  x_421 & ~n_20365;
assign n_20367 = ~x_421 &  n_20365;
assign n_20368 = ~n_20366 & ~n_20367;
assign n_20369 =  x_420 & ~n_20332;
assign n_20370 =  x_100 &  n_20332;
assign n_20371 = ~n_20369 & ~n_20370;
assign n_20372 =  x_420 & ~n_20371;
assign n_20373 = ~x_420 &  n_20371;
assign n_20374 = ~n_20372 & ~n_20373;
assign n_20375 =  x_419 & ~n_20332;
assign n_20376 =  x_99 &  n_20332;
assign n_20377 = ~n_20375 & ~n_20376;
assign n_20378 =  x_419 & ~n_20377;
assign n_20379 = ~x_419 &  n_20377;
assign n_20380 = ~n_20378 & ~n_20379;
assign n_20381 =  x_418 & ~n_20332;
assign n_20382 =  x_98 &  n_20332;
assign n_20383 = ~n_20381 & ~n_20382;
assign n_20384 =  x_418 & ~n_20383;
assign n_20385 = ~x_418 &  n_20383;
assign n_20386 = ~n_20384 & ~n_20385;
assign n_20387 =  x_417 & ~n_20332;
assign n_20388 =  x_97 &  n_20332;
assign n_20389 = ~n_20387 & ~n_20388;
assign n_20390 =  x_417 & ~n_20389;
assign n_20391 = ~x_417 &  n_20389;
assign n_20392 = ~n_20390 & ~n_20391;
assign n_20393 =  x_416 & ~n_20332;
assign n_20394 =  x_96 &  n_20332;
assign n_20395 = ~n_20393 & ~n_20394;
assign n_20396 =  x_416 & ~n_20395;
assign n_20397 = ~x_416 &  n_20395;
assign n_20398 = ~n_20396 & ~n_20397;
assign n_20399 =  x_415 & ~n_20332;
assign n_20400 =  x_95 &  n_20332;
assign n_20401 = ~n_20399 & ~n_20400;
assign n_20402 =  x_415 & ~n_20401;
assign n_20403 = ~x_415 &  n_20401;
assign n_20404 = ~n_20402 & ~n_20403;
assign n_20405 =  x_414 & ~n_20332;
assign n_20406 =  x_94 &  n_20332;
assign n_20407 = ~n_20405 & ~n_20406;
assign n_20408 =  x_414 & ~n_20407;
assign n_20409 = ~x_414 &  n_20407;
assign n_20410 = ~n_20408 & ~n_20409;
assign n_20411 =  x_413 & ~n_20332;
assign n_20412 =  x_93 &  n_20332;
assign n_20413 = ~n_20411 & ~n_20412;
assign n_20414 =  x_413 & ~n_20413;
assign n_20415 = ~x_413 &  n_20413;
assign n_20416 = ~n_20414 & ~n_20415;
assign n_20417 =  x_412 & ~n_20332;
assign n_20418 =  x_92 &  n_20332;
assign n_20419 = ~n_20417 & ~n_20418;
assign n_20420 =  x_412 & ~n_20419;
assign n_20421 = ~x_412 &  n_20419;
assign n_20422 = ~n_20420 & ~n_20421;
assign n_20423 =  x_411 & ~n_20332;
assign n_20424 =  x_91 &  n_20332;
assign n_20425 = ~n_20423 & ~n_20424;
assign n_20426 =  x_411 & ~n_20425;
assign n_20427 = ~x_411 &  n_20425;
assign n_20428 = ~n_20426 & ~n_20427;
assign n_20429 =  x_410 & ~n_20332;
assign n_20430 =  x_90 &  n_20332;
assign n_20431 = ~n_20429 & ~n_20430;
assign n_20432 =  x_410 & ~n_20431;
assign n_20433 = ~x_410 &  n_20431;
assign n_20434 = ~n_20432 & ~n_20433;
assign n_20435 =  x_409 & ~n_20332;
assign n_20436 =  x_89 &  n_20332;
assign n_20437 = ~n_20435 & ~n_20436;
assign n_20438 =  x_409 & ~n_20437;
assign n_20439 = ~x_409 &  n_20437;
assign n_20440 = ~n_20438 & ~n_20439;
assign n_20441 =  x_408 & ~n_20332;
assign n_20442 =  x_88 &  n_20332;
assign n_20443 = ~n_20441 & ~n_20442;
assign n_20444 =  x_408 & ~n_20443;
assign n_20445 = ~x_408 &  n_20443;
assign n_20446 = ~n_20444 & ~n_20445;
assign n_20447 =  x_407 & ~n_20332;
assign n_20448 =  x_87 &  n_20332;
assign n_20449 = ~n_20447 & ~n_20448;
assign n_20450 =  x_407 & ~n_20449;
assign n_20451 = ~x_407 &  n_20449;
assign n_20452 = ~n_20450 & ~n_20451;
assign n_20453 =  x_406 & ~n_20332;
assign n_20454 =  x_86 &  n_20332;
assign n_20455 = ~n_20453 & ~n_20454;
assign n_20456 =  x_406 & ~n_20455;
assign n_20457 = ~x_406 &  n_20455;
assign n_20458 = ~n_20456 & ~n_20457;
assign n_20459 =  x_405 & ~n_20332;
assign n_20460 =  x_85 &  n_20332;
assign n_20461 = ~n_20459 & ~n_20460;
assign n_20462 =  x_405 & ~n_20461;
assign n_20463 = ~x_405 &  n_20461;
assign n_20464 = ~n_20462 & ~n_20463;
assign n_20465 =  x_404 & ~n_20332;
assign n_20466 =  x_84 &  n_20332;
assign n_20467 = ~n_20465 & ~n_20466;
assign n_20468 =  x_404 & ~n_20467;
assign n_20469 = ~x_404 &  n_20467;
assign n_20470 = ~n_20468 & ~n_20469;
assign n_20471 =  x_403 & ~n_20332;
assign n_20472 =  x_83 &  n_20332;
assign n_20473 = ~n_20471 & ~n_20472;
assign n_20474 =  x_403 & ~n_20473;
assign n_20475 = ~x_403 &  n_20473;
assign n_20476 = ~n_20474 & ~n_20475;
assign n_20477 =  x_402 & ~n_20332;
assign n_20478 =  x_82 &  n_20332;
assign n_20479 = ~n_20477 & ~n_20478;
assign n_20480 =  x_402 & ~n_20479;
assign n_20481 = ~x_402 &  n_20479;
assign n_20482 = ~n_20480 & ~n_20481;
assign n_20483 =  x_401 & ~n_20332;
assign n_20484 =  x_81 &  n_20332;
assign n_20485 = ~n_20483 & ~n_20484;
assign n_20486 =  x_401 & ~n_20485;
assign n_20487 = ~x_401 &  n_20485;
assign n_20488 = ~n_20486 & ~n_20487;
assign n_20489 =  x_400 & ~n_20332;
assign n_20490 =  x_80 &  n_20332;
assign n_20491 = ~n_20489 & ~n_20490;
assign n_20492 =  x_400 & ~n_20491;
assign n_20493 = ~x_400 &  n_20491;
assign n_20494 = ~n_20492 & ~n_20493;
assign n_20495 =  x_399 & ~n_20332;
assign n_20496 =  x_79 &  n_20332;
assign n_20497 = ~n_20495 & ~n_20496;
assign n_20498 =  x_399 & ~n_20497;
assign n_20499 = ~x_399 &  n_20497;
assign n_20500 = ~n_20498 & ~n_20499;
assign n_20501 =  x_398 & ~n_20332;
assign n_20502 =  x_78 &  n_20332;
assign n_20503 = ~n_20501 & ~n_20502;
assign n_20504 =  x_398 & ~n_20503;
assign n_20505 = ~x_398 &  n_20503;
assign n_20506 = ~n_20504 & ~n_20505;
assign n_20507 =  x_397 & ~n_20332;
assign n_20508 =  x_77 &  n_20332;
assign n_20509 = ~n_20507 & ~n_20508;
assign n_20510 =  x_397 & ~n_20509;
assign n_20511 = ~x_397 &  n_20509;
assign n_20512 = ~n_20510 & ~n_20511;
assign n_20513 =  x_396 & ~n_20332;
assign n_20514 =  x_76 &  n_20332;
assign n_20515 = ~n_20513 & ~n_20514;
assign n_20516 =  x_396 & ~n_20515;
assign n_20517 = ~x_396 &  n_20515;
assign n_20518 = ~n_20516 & ~n_20517;
assign n_20519 =  x_395 & ~n_20332;
assign n_20520 =  x_75 &  n_20332;
assign n_20521 = ~n_20519 & ~n_20520;
assign n_20522 =  x_395 & ~n_20521;
assign n_20523 = ~x_395 &  n_20521;
assign n_20524 = ~n_20522 & ~n_20523;
assign n_20525 =  n_1906 &  n_18439;
assign n_20526 =  x_394 & ~n_20525;
assign n_20527 =  i_32 &  n_20525;
assign n_20528 = ~n_20526 & ~n_20527;
assign n_20529 =  x_394 & ~n_20528;
assign n_20530 = ~x_394 &  n_20528;
assign n_20531 = ~n_20529 & ~n_20530;
assign n_20532 =  x_393 & ~n_20525;
assign n_20533 =  i_31 &  n_20525;
assign n_20534 = ~n_20532 & ~n_20533;
assign n_20535 =  x_393 & ~n_20534;
assign n_20536 = ~x_393 &  n_20534;
assign n_20537 = ~n_20535 & ~n_20536;
assign n_20538 =  x_392 & ~n_20525;
assign n_20539 =  i_30 &  n_20525;
assign n_20540 = ~n_20538 & ~n_20539;
assign n_20541 =  x_392 & ~n_20540;
assign n_20542 = ~x_392 &  n_20540;
assign n_20543 = ~n_20541 & ~n_20542;
assign n_20544 =  x_391 & ~n_20525;
assign n_20545 =  i_29 &  n_20525;
assign n_20546 = ~n_20544 & ~n_20545;
assign n_20547 =  x_391 & ~n_20546;
assign n_20548 = ~x_391 &  n_20546;
assign n_20549 = ~n_20547 & ~n_20548;
assign n_20550 =  x_390 & ~n_20525;
assign n_20551 =  i_28 &  n_20525;
assign n_20552 = ~n_20550 & ~n_20551;
assign n_20553 =  x_390 & ~n_20552;
assign n_20554 = ~x_390 &  n_20552;
assign n_20555 = ~n_20553 & ~n_20554;
assign n_20556 =  x_389 & ~n_20525;
assign n_20557 =  i_27 &  n_20525;
assign n_20558 = ~n_20556 & ~n_20557;
assign n_20559 =  x_389 & ~n_20558;
assign n_20560 = ~x_389 &  n_20558;
assign n_20561 = ~n_20559 & ~n_20560;
assign n_20562 =  x_388 & ~n_20525;
assign n_20563 =  i_26 &  n_20525;
assign n_20564 = ~n_20562 & ~n_20563;
assign n_20565 =  x_388 & ~n_20564;
assign n_20566 = ~x_388 &  n_20564;
assign n_20567 = ~n_20565 & ~n_20566;
assign n_20568 =  x_387 & ~n_20525;
assign n_20569 =  i_25 &  n_20525;
assign n_20570 = ~n_20568 & ~n_20569;
assign n_20571 =  x_387 & ~n_20570;
assign n_20572 = ~x_387 &  n_20570;
assign n_20573 = ~n_20571 & ~n_20572;
assign n_20574 =  x_386 & ~n_20525;
assign n_20575 =  i_24 &  n_20525;
assign n_20576 = ~n_20574 & ~n_20575;
assign n_20577 =  x_386 & ~n_20576;
assign n_20578 = ~x_386 &  n_20576;
assign n_20579 = ~n_20577 & ~n_20578;
assign n_20580 =  x_385 & ~n_20525;
assign n_20581 =  i_23 &  n_20525;
assign n_20582 = ~n_20580 & ~n_20581;
assign n_20583 =  x_385 & ~n_20582;
assign n_20584 = ~x_385 &  n_20582;
assign n_20585 = ~n_20583 & ~n_20584;
assign n_20586 =  x_384 & ~n_20525;
assign n_20587 =  i_22 &  n_20525;
assign n_20588 = ~n_20586 & ~n_20587;
assign n_20589 =  x_384 & ~n_20588;
assign n_20590 = ~x_384 &  n_20588;
assign n_20591 = ~n_20589 & ~n_20590;
assign n_20592 =  x_383 & ~n_20525;
assign n_20593 =  i_21 &  n_20525;
assign n_20594 = ~n_20592 & ~n_20593;
assign n_20595 =  x_383 & ~n_20594;
assign n_20596 = ~x_383 &  n_20594;
assign n_20597 = ~n_20595 & ~n_20596;
assign n_20598 =  x_382 & ~n_20525;
assign n_20599 =  i_20 &  n_20525;
assign n_20600 = ~n_20598 & ~n_20599;
assign n_20601 =  x_382 & ~n_20600;
assign n_20602 = ~x_382 &  n_20600;
assign n_20603 = ~n_20601 & ~n_20602;
assign n_20604 =  x_381 & ~n_20525;
assign n_20605 =  i_19 &  n_20525;
assign n_20606 = ~n_20604 & ~n_20605;
assign n_20607 =  x_381 & ~n_20606;
assign n_20608 = ~x_381 &  n_20606;
assign n_20609 = ~n_20607 & ~n_20608;
assign n_20610 =  x_380 & ~n_20525;
assign n_20611 =  i_18 &  n_20525;
assign n_20612 = ~n_20610 & ~n_20611;
assign n_20613 =  x_380 & ~n_20612;
assign n_20614 = ~x_380 &  n_20612;
assign n_20615 = ~n_20613 & ~n_20614;
assign n_20616 =  x_379 & ~n_20525;
assign n_20617 =  i_17 &  n_20525;
assign n_20618 = ~n_20616 & ~n_20617;
assign n_20619 =  x_379 & ~n_20618;
assign n_20620 = ~x_379 &  n_20618;
assign n_20621 = ~n_20619 & ~n_20620;
assign n_20622 =  x_378 & ~n_20525;
assign n_20623 =  i_16 &  n_20525;
assign n_20624 = ~n_20622 & ~n_20623;
assign n_20625 =  x_378 & ~n_20624;
assign n_20626 = ~x_378 &  n_20624;
assign n_20627 = ~n_20625 & ~n_20626;
assign n_20628 =  x_377 & ~n_20525;
assign n_20629 =  i_15 &  n_20525;
assign n_20630 = ~n_20628 & ~n_20629;
assign n_20631 =  x_377 & ~n_20630;
assign n_20632 = ~x_377 &  n_20630;
assign n_20633 = ~n_20631 & ~n_20632;
assign n_20634 =  x_376 & ~n_20525;
assign n_20635 =  i_14 &  n_20525;
assign n_20636 = ~n_20634 & ~n_20635;
assign n_20637 =  x_376 & ~n_20636;
assign n_20638 = ~x_376 &  n_20636;
assign n_20639 = ~n_20637 & ~n_20638;
assign n_20640 =  x_375 & ~n_20525;
assign n_20641 =  i_13 &  n_20525;
assign n_20642 = ~n_20640 & ~n_20641;
assign n_20643 =  x_375 & ~n_20642;
assign n_20644 = ~x_375 &  n_20642;
assign n_20645 = ~n_20643 & ~n_20644;
assign n_20646 =  x_374 & ~n_20525;
assign n_20647 =  i_12 &  n_20525;
assign n_20648 = ~n_20646 & ~n_20647;
assign n_20649 =  x_374 & ~n_20648;
assign n_20650 = ~x_374 &  n_20648;
assign n_20651 = ~n_20649 & ~n_20650;
assign n_20652 =  x_373 & ~n_20525;
assign n_20653 =  i_11 &  n_20525;
assign n_20654 = ~n_20652 & ~n_20653;
assign n_20655 =  x_373 & ~n_20654;
assign n_20656 = ~x_373 &  n_20654;
assign n_20657 = ~n_20655 & ~n_20656;
assign n_20658 =  x_372 & ~n_20525;
assign n_20659 =  i_10 &  n_20525;
assign n_20660 = ~n_20658 & ~n_20659;
assign n_20661 =  x_372 & ~n_20660;
assign n_20662 = ~x_372 &  n_20660;
assign n_20663 = ~n_20661 & ~n_20662;
assign n_20664 =  x_371 & ~n_20525;
assign n_20665 =  i_9 &  n_20525;
assign n_20666 = ~n_20664 & ~n_20665;
assign n_20667 =  x_371 & ~n_20666;
assign n_20668 = ~x_371 &  n_20666;
assign n_20669 = ~n_20667 & ~n_20668;
assign n_20670 =  x_370 & ~n_20525;
assign n_20671 =  i_8 &  n_20525;
assign n_20672 = ~n_20670 & ~n_20671;
assign n_20673 =  x_370 & ~n_20672;
assign n_20674 = ~x_370 &  n_20672;
assign n_20675 = ~n_20673 & ~n_20674;
assign n_20676 =  x_369 & ~n_20525;
assign n_20677 =  i_7 &  n_20525;
assign n_20678 = ~n_20676 & ~n_20677;
assign n_20679 =  x_369 & ~n_20678;
assign n_20680 = ~x_369 &  n_20678;
assign n_20681 = ~n_20679 & ~n_20680;
assign n_20682 =  x_368 & ~n_20525;
assign n_20683 =  i_6 &  n_20525;
assign n_20684 = ~n_20682 & ~n_20683;
assign n_20685 =  x_368 & ~n_20684;
assign n_20686 = ~x_368 &  n_20684;
assign n_20687 = ~n_20685 & ~n_20686;
assign n_20688 =  x_367 & ~n_20525;
assign n_20689 =  i_5 &  n_20525;
assign n_20690 = ~n_20688 & ~n_20689;
assign n_20691 =  x_367 & ~n_20690;
assign n_20692 = ~x_367 &  n_20690;
assign n_20693 = ~n_20691 & ~n_20692;
assign n_20694 =  x_366 & ~n_20525;
assign n_20695 =  i_4 &  n_20525;
assign n_20696 = ~n_20694 & ~n_20695;
assign n_20697 =  x_366 & ~n_20696;
assign n_20698 = ~x_366 &  n_20696;
assign n_20699 = ~n_20697 & ~n_20698;
assign n_20700 =  x_365 & ~n_20525;
assign n_20701 =  i_3 &  n_20525;
assign n_20702 = ~n_20700 & ~n_20701;
assign n_20703 =  x_365 & ~n_20702;
assign n_20704 = ~x_365 &  n_20702;
assign n_20705 = ~n_20703 & ~n_20704;
assign n_20706 =  x_364 & ~n_20525;
assign n_20707 =  i_2 &  n_20525;
assign n_20708 = ~n_20706 & ~n_20707;
assign n_20709 =  x_364 & ~n_20708;
assign n_20710 = ~x_364 &  n_20708;
assign n_20711 = ~n_20709 & ~n_20710;
assign n_20712 =  x_363 & ~n_20525;
assign n_20713 =  i_1 &  n_20525;
assign n_20714 = ~n_20712 & ~n_20713;
assign n_20715 =  x_363 & ~n_20714;
assign n_20716 = ~x_363 &  n_20714;
assign n_20717 = ~n_20715 & ~n_20716;
assign n_20718 =  n_1314 &  n_6332;
assign n_20719 =  n_8059 &  n_7865;
assign n_20720 = ~n_20718 & ~n_20719;
assign n_20721 =  x_42 & ~n_20720;
assign n_20722 =  x_362 & ~n_20721;
assign n_20723 =  i_32 &  n_20721;
assign n_20724 = ~n_20722 & ~n_20723;
assign n_20725 =  x_362 & ~n_20724;
assign n_20726 = ~x_362 &  n_20724;
assign n_20727 = ~n_20725 & ~n_20726;
assign n_20728 =  x_361 & ~n_20721;
assign n_20729 =  i_31 &  n_20721;
assign n_20730 = ~n_20728 & ~n_20729;
assign n_20731 =  x_361 & ~n_20730;
assign n_20732 = ~x_361 &  n_20730;
assign n_20733 = ~n_20731 & ~n_20732;
assign n_20734 =  x_360 & ~n_20721;
assign n_20735 =  i_30 &  n_20721;
assign n_20736 = ~n_20734 & ~n_20735;
assign n_20737 =  x_360 & ~n_20736;
assign n_20738 = ~x_360 &  n_20736;
assign n_20739 = ~n_20737 & ~n_20738;
assign n_20740 =  x_359 & ~n_20721;
assign n_20741 =  i_29 &  n_20721;
assign n_20742 = ~n_20740 & ~n_20741;
assign n_20743 =  x_359 & ~n_20742;
assign n_20744 = ~x_359 &  n_20742;
assign n_20745 = ~n_20743 & ~n_20744;
assign n_20746 =  x_358 & ~n_20721;
assign n_20747 =  i_28 &  n_20721;
assign n_20748 = ~n_20746 & ~n_20747;
assign n_20749 =  x_358 & ~n_20748;
assign n_20750 = ~x_358 &  n_20748;
assign n_20751 = ~n_20749 & ~n_20750;
assign n_20752 =  x_357 & ~n_20721;
assign n_20753 =  i_27 &  n_20721;
assign n_20754 = ~n_20752 & ~n_20753;
assign n_20755 =  x_357 & ~n_20754;
assign n_20756 = ~x_357 &  n_20754;
assign n_20757 = ~n_20755 & ~n_20756;
assign n_20758 =  x_356 & ~n_20721;
assign n_20759 =  i_26 &  n_20721;
assign n_20760 = ~n_20758 & ~n_20759;
assign n_20761 =  x_356 & ~n_20760;
assign n_20762 = ~x_356 &  n_20760;
assign n_20763 = ~n_20761 & ~n_20762;
assign n_20764 =  x_355 & ~n_20721;
assign n_20765 =  i_25 &  n_20721;
assign n_20766 = ~n_20764 & ~n_20765;
assign n_20767 =  x_355 & ~n_20766;
assign n_20768 = ~x_355 &  n_20766;
assign n_20769 = ~n_20767 & ~n_20768;
assign n_20770 =  x_354 & ~n_20721;
assign n_20771 =  i_24 &  n_20721;
assign n_20772 = ~n_20770 & ~n_20771;
assign n_20773 =  x_354 & ~n_20772;
assign n_20774 = ~x_354 &  n_20772;
assign n_20775 = ~n_20773 & ~n_20774;
assign n_20776 =  x_353 & ~n_20721;
assign n_20777 =  i_23 &  n_20721;
assign n_20778 = ~n_20776 & ~n_20777;
assign n_20779 =  x_353 & ~n_20778;
assign n_20780 = ~x_353 &  n_20778;
assign n_20781 = ~n_20779 & ~n_20780;
assign n_20782 =  x_352 & ~n_20721;
assign n_20783 =  i_22 &  n_20721;
assign n_20784 = ~n_20782 & ~n_20783;
assign n_20785 =  x_352 & ~n_20784;
assign n_20786 = ~x_352 &  n_20784;
assign n_20787 = ~n_20785 & ~n_20786;
assign n_20788 =  x_351 & ~n_20721;
assign n_20789 =  i_21 &  n_20721;
assign n_20790 = ~n_20788 & ~n_20789;
assign n_20791 =  x_351 & ~n_20790;
assign n_20792 = ~x_351 &  n_20790;
assign n_20793 = ~n_20791 & ~n_20792;
assign n_20794 =  x_350 & ~n_20721;
assign n_20795 =  i_20 &  n_20721;
assign n_20796 = ~n_20794 & ~n_20795;
assign n_20797 =  x_350 & ~n_20796;
assign n_20798 = ~x_350 &  n_20796;
assign n_20799 = ~n_20797 & ~n_20798;
assign n_20800 =  x_349 & ~n_20721;
assign n_20801 =  i_19 &  n_20721;
assign n_20802 = ~n_20800 & ~n_20801;
assign n_20803 =  x_349 & ~n_20802;
assign n_20804 = ~x_349 &  n_20802;
assign n_20805 = ~n_20803 & ~n_20804;
assign n_20806 =  x_348 & ~n_20721;
assign n_20807 =  i_18 &  n_20721;
assign n_20808 = ~n_20806 & ~n_20807;
assign n_20809 =  x_348 & ~n_20808;
assign n_20810 = ~x_348 &  n_20808;
assign n_20811 = ~n_20809 & ~n_20810;
assign n_20812 =  x_347 & ~n_20721;
assign n_20813 =  i_17 &  n_20721;
assign n_20814 = ~n_20812 & ~n_20813;
assign n_20815 =  x_347 & ~n_20814;
assign n_20816 = ~x_347 &  n_20814;
assign n_20817 = ~n_20815 & ~n_20816;
assign n_20818 =  x_346 & ~n_20721;
assign n_20819 =  i_16 &  n_20721;
assign n_20820 = ~n_20818 & ~n_20819;
assign n_20821 =  x_346 & ~n_20820;
assign n_20822 = ~x_346 &  n_20820;
assign n_20823 = ~n_20821 & ~n_20822;
assign n_20824 =  x_345 & ~n_20721;
assign n_20825 =  i_15 &  n_20721;
assign n_20826 = ~n_20824 & ~n_20825;
assign n_20827 =  x_345 & ~n_20826;
assign n_20828 = ~x_345 &  n_20826;
assign n_20829 = ~n_20827 & ~n_20828;
assign n_20830 =  x_344 & ~n_20721;
assign n_20831 =  i_14 &  n_20721;
assign n_20832 = ~n_20830 & ~n_20831;
assign n_20833 =  x_344 & ~n_20832;
assign n_20834 = ~x_344 &  n_20832;
assign n_20835 = ~n_20833 & ~n_20834;
assign n_20836 =  x_343 & ~n_20721;
assign n_20837 =  i_13 &  n_20721;
assign n_20838 = ~n_20836 & ~n_20837;
assign n_20839 =  x_343 & ~n_20838;
assign n_20840 = ~x_343 &  n_20838;
assign n_20841 = ~n_20839 & ~n_20840;
assign n_20842 =  x_342 & ~n_20721;
assign n_20843 =  i_12 &  n_20721;
assign n_20844 = ~n_20842 & ~n_20843;
assign n_20845 =  x_342 & ~n_20844;
assign n_20846 = ~x_342 &  n_20844;
assign n_20847 = ~n_20845 & ~n_20846;
assign n_20848 =  x_341 & ~n_20721;
assign n_20849 =  i_11 &  n_20721;
assign n_20850 = ~n_20848 & ~n_20849;
assign n_20851 =  x_341 & ~n_20850;
assign n_20852 = ~x_341 &  n_20850;
assign n_20853 = ~n_20851 & ~n_20852;
assign n_20854 =  x_340 & ~n_20721;
assign n_20855 =  i_10 &  n_20721;
assign n_20856 = ~n_20854 & ~n_20855;
assign n_20857 =  x_340 & ~n_20856;
assign n_20858 = ~x_340 &  n_20856;
assign n_20859 = ~n_20857 & ~n_20858;
assign n_20860 =  x_339 & ~n_20721;
assign n_20861 =  i_9 &  n_20721;
assign n_20862 = ~n_20860 & ~n_20861;
assign n_20863 =  x_339 & ~n_20862;
assign n_20864 = ~x_339 &  n_20862;
assign n_20865 = ~n_20863 & ~n_20864;
assign n_20866 =  x_338 & ~n_20721;
assign n_20867 =  i_8 &  n_20721;
assign n_20868 = ~n_20866 & ~n_20867;
assign n_20869 =  x_338 & ~n_20868;
assign n_20870 = ~x_338 &  n_20868;
assign n_20871 = ~n_20869 & ~n_20870;
assign n_20872 =  x_337 & ~n_20721;
assign n_20873 =  i_7 &  n_20721;
assign n_20874 = ~n_20872 & ~n_20873;
assign n_20875 =  x_337 & ~n_20874;
assign n_20876 = ~x_337 &  n_20874;
assign n_20877 = ~n_20875 & ~n_20876;
assign n_20878 =  x_336 & ~n_20721;
assign n_20879 =  i_6 &  n_20721;
assign n_20880 = ~n_20878 & ~n_20879;
assign n_20881 =  x_336 & ~n_20880;
assign n_20882 = ~x_336 &  n_20880;
assign n_20883 = ~n_20881 & ~n_20882;
assign n_20884 =  x_335 & ~n_20721;
assign n_20885 =  i_5 &  n_20721;
assign n_20886 = ~n_20884 & ~n_20885;
assign n_20887 =  x_335 & ~n_20886;
assign n_20888 = ~x_335 &  n_20886;
assign n_20889 = ~n_20887 & ~n_20888;
assign n_20890 =  x_334 & ~n_20721;
assign n_20891 =  i_4 &  n_20721;
assign n_20892 = ~n_20890 & ~n_20891;
assign n_20893 =  x_334 & ~n_20892;
assign n_20894 = ~x_334 &  n_20892;
assign n_20895 = ~n_20893 & ~n_20894;
assign n_20896 =  x_333 & ~n_20721;
assign n_20897 =  i_3 &  n_20721;
assign n_20898 = ~n_20896 & ~n_20897;
assign n_20899 =  x_333 & ~n_20898;
assign n_20900 = ~x_333 &  n_20898;
assign n_20901 = ~n_20899 & ~n_20900;
assign n_20902 =  x_332 & ~n_20721;
assign n_20903 =  i_2 &  n_20721;
assign n_20904 = ~n_20902 & ~n_20903;
assign n_20905 =  x_332 & ~n_20904;
assign n_20906 = ~x_332 &  n_20904;
assign n_20907 = ~n_20905 & ~n_20906;
assign n_20908 =  x_331 & ~n_20721;
assign n_20909 =  i_1 &  n_20721;
assign n_20910 = ~n_20908 & ~n_20909;
assign n_20911 =  x_331 & ~n_20910;
assign n_20912 = ~x_331 &  n_20910;
assign n_20913 = ~n_20911 & ~n_20912;
assign n_20914 =  n_8818 &  n_18439;
assign n_20915 =  x_330 & ~n_20914;
assign n_20916 =  i_32 &  n_20914;
assign n_20917 = ~n_20915 & ~n_20916;
assign n_20918 =  x_330 & ~n_20917;
assign n_20919 = ~x_330 &  n_20917;
assign n_20920 = ~n_20918 & ~n_20919;
assign n_20921 =  x_329 & ~n_20914;
assign n_20922 =  i_31 &  n_20914;
assign n_20923 = ~n_20921 & ~n_20922;
assign n_20924 =  x_329 & ~n_20923;
assign n_20925 = ~x_329 &  n_20923;
assign n_20926 = ~n_20924 & ~n_20925;
assign n_20927 =  x_328 & ~n_20914;
assign n_20928 =  i_30 &  n_20914;
assign n_20929 = ~n_20927 & ~n_20928;
assign n_20930 =  x_328 & ~n_20929;
assign n_20931 = ~x_328 &  n_20929;
assign n_20932 = ~n_20930 & ~n_20931;
assign n_20933 =  x_327 & ~n_20914;
assign n_20934 =  i_29 &  n_20914;
assign n_20935 = ~n_20933 & ~n_20934;
assign n_20936 =  x_327 & ~n_20935;
assign n_20937 = ~x_327 &  n_20935;
assign n_20938 = ~n_20936 & ~n_20937;
assign n_20939 =  x_326 & ~n_20914;
assign n_20940 =  i_28 &  n_20914;
assign n_20941 = ~n_20939 & ~n_20940;
assign n_20942 =  x_326 & ~n_20941;
assign n_20943 = ~x_326 &  n_20941;
assign n_20944 = ~n_20942 & ~n_20943;
assign n_20945 =  x_325 & ~n_20914;
assign n_20946 =  i_27 &  n_20914;
assign n_20947 = ~n_20945 & ~n_20946;
assign n_20948 =  x_325 & ~n_20947;
assign n_20949 = ~x_325 &  n_20947;
assign n_20950 = ~n_20948 & ~n_20949;
assign n_20951 =  x_324 & ~n_20914;
assign n_20952 =  i_26 &  n_20914;
assign n_20953 = ~n_20951 & ~n_20952;
assign n_20954 =  x_324 & ~n_20953;
assign n_20955 = ~x_324 &  n_20953;
assign n_20956 = ~n_20954 & ~n_20955;
assign n_20957 =  x_323 & ~n_20914;
assign n_20958 =  i_25 &  n_20914;
assign n_20959 = ~n_20957 & ~n_20958;
assign n_20960 =  x_323 & ~n_20959;
assign n_20961 = ~x_323 &  n_20959;
assign n_20962 = ~n_20960 & ~n_20961;
assign n_20963 =  x_322 & ~n_20914;
assign n_20964 =  i_24 &  n_20914;
assign n_20965 = ~n_20963 & ~n_20964;
assign n_20966 =  x_322 & ~n_20965;
assign n_20967 = ~x_322 &  n_20965;
assign n_20968 = ~n_20966 & ~n_20967;
assign n_20969 =  x_321 & ~n_20914;
assign n_20970 =  i_23 &  n_20914;
assign n_20971 = ~n_20969 & ~n_20970;
assign n_20972 =  x_321 & ~n_20971;
assign n_20973 = ~x_321 &  n_20971;
assign n_20974 = ~n_20972 & ~n_20973;
assign n_20975 =  x_320 & ~n_20914;
assign n_20976 =  i_22 &  n_20914;
assign n_20977 = ~n_20975 & ~n_20976;
assign n_20978 =  x_320 & ~n_20977;
assign n_20979 = ~x_320 &  n_20977;
assign n_20980 = ~n_20978 & ~n_20979;
assign n_20981 =  x_319 & ~n_20914;
assign n_20982 =  i_21 &  n_20914;
assign n_20983 = ~n_20981 & ~n_20982;
assign n_20984 =  x_319 & ~n_20983;
assign n_20985 = ~x_319 &  n_20983;
assign n_20986 = ~n_20984 & ~n_20985;
assign n_20987 =  x_318 & ~n_20914;
assign n_20988 =  i_20 &  n_20914;
assign n_20989 = ~n_20987 & ~n_20988;
assign n_20990 =  x_318 & ~n_20989;
assign n_20991 = ~x_318 &  n_20989;
assign n_20992 = ~n_20990 & ~n_20991;
assign n_20993 =  x_317 & ~n_20914;
assign n_20994 =  i_19 &  n_20914;
assign n_20995 = ~n_20993 & ~n_20994;
assign n_20996 =  x_317 & ~n_20995;
assign n_20997 = ~x_317 &  n_20995;
assign n_20998 = ~n_20996 & ~n_20997;
assign n_20999 =  x_316 & ~n_20914;
assign n_21000 =  i_18 &  n_20914;
assign n_21001 = ~n_20999 & ~n_21000;
assign n_21002 =  x_316 & ~n_21001;
assign n_21003 = ~x_316 &  n_21001;
assign n_21004 = ~n_21002 & ~n_21003;
assign n_21005 =  x_315 & ~n_20914;
assign n_21006 =  i_17 &  n_20914;
assign n_21007 = ~n_21005 & ~n_21006;
assign n_21008 =  x_315 & ~n_21007;
assign n_21009 = ~x_315 &  n_21007;
assign n_21010 = ~n_21008 & ~n_21009;
assign n_21011 =  x_314 & ~n_20914;
assign n_21012 =  i_16 &  n_20914;
assign n_21013 = ~n_21011 & ~n_21012;
assign n_21014 =  x_314 & ~n_21013;
assign n_21015 = ~x_314 &  n_21013;
assign n_21016 = ~n_21014 & ~n_21015;
assign n_21017 =  x_313 & ~n_20914;
assign n_21018 =  i_15 &  n_20914;
assign n_21019 = ~n_21017 & ~n_21018;
assign n_21020 =  x_313 & ~n_21019;
assign n_21021 = ~x_313 &  n_21019;
assign n_21022 = ~n_21020 & ~n_21021;
assign n_21023 =  x_312 & ~n_20914;
assign n_21024 =  i_14 &  n_20914;
assign n_21025 = ~n_21023 & ~n_21024;
assign n_21026 =  x_312 & ~n_21025;
assign n_21027 = ~x_312 &  n_21025;
assign n_21028 = ~n_21026 & ~n_21027;
assign n_21029 =  x_311 & ~n_20914;
assign n_21030 =  i_13 &  n_20914;
assign n_21031 = ~n_21029 & ~n_21030;
assign n_21032 =  x_311 & ~n_21031;
assign n_21033 = ~x_311 &  n_21031;
assign n_21034 = ~n_21032 & ~n_21033;
assign n_21035 =  x_310 & ~n_20914;
assign n_21036 =  i_12 &  n_20914;
assign n_21037 = ~n_21035 & ~n_21036;
assign n_21038 =  x_310 & ~n_21037;
assign n_21039 = ~x_310 &  n_21037;
assign n_21040 = ~n_21038 & ~n_21039;
assign n_21041 =  x_309 & ~n_20914;
assign n_21042 =  i_11 &  n_20914;
assign n_21043 = ~n_21041 & ~n_21042;
assign n_21044 =  x_309 & ~n_21043;
assign n_21045 = ~x_309 &  n_21043;
assign n_21046 = ~n_21044 & ~n_21045;
assign n_21047 =  x_308 & ~n_20914;
assign n_21048 =  i_10 &  n_20914;
assign n_21049 = ~n_21047 & ~n_21048;
assign n_21050 =  x_308 & ~n_21049;
assign n_21051 = ~x_308 &  n_21049;
assign n_21052 = ~n_21050 & ~n_21051;
assign n_21053 =  x_307 & ~n_20914;
assign n_21054 =  i_9 &  n_20914;
assign n_21055 = ~n_21053 & ~n_21054;
assign n_21056 =  x_307 & ~n_21055;
assign n_21057 = ~x_307 &  n_21055;
assign n_21058 = ~n_21056 & ~n_21057;
assign n_21059 =  x_306 & ~n_20914;
assign n_21060 =  i_8 &  n_20914;
assign n_21061 = ~n_21059 & ~n_21060;
assign n_21062 =  x_306 & ~n_21061;
assign n_21063 = ~x_306 &  n_21061;
assign n_21064 = ~n_21062 & ~n_21063;
assign n_21065 =  x_305 & ~n_20914;
assign n_21066 =  i_7 &  n_20914;
assign n_21067 = ~n_21065 & ~n_21066;
assign n_21068 =  x_305 & ~n_21067;
assign n_21069 = ~x_305 &  n_21067;
assign n_21070 = ~n_21068 & ~n_21069;
assign n_21071 =  x_304 & ~n_20914;
assign n_21072 =  i_6 &  n_20914;
assign n_21073 = ~n_21071 & ~n_21072;
assign n_21074 =  x_304 & ~n_21073;
assign n_21075 = ~x_304 &  n_21073;
assign n_21076 = ~n_21074 & ~n_21075;
assign n_21077 =  x_303 & ~n_20914;
assign n_21078 =  i_5 &  n_20914;
assign n_21079 = ~n_21077 & ~n_21078;
assign n_21080 =  x_303 & ~n_21079;
assign n_21081 = ~x_303 &  n_21079;
assign n_21082 = ~n_21080 & ~n_21081;
assign n_21083 =  x_302 & ~n_20914;
assign n_21084 =  i_4 &  n_20914;
assign n_21085 = ~n_21083 & ~n_21084;
assign n_21086 =  x_302 & ~n_21085;
assign n_21087 = ~x_302 &  n_21085;
assign n_21088 = ~n_21086 & ~n_21087;
assign n_21089 =  x_301 & ~n_20914;
assign n_21090 =  i_3 &  n_20914;
assign n_21091 = ~n_21089 & ~n_21090;
assign n_21092 =  x_301 & ~n_21091;
assign n_21093 = ~x_301 &  n_21091;
assign n_21094 = ~n_21092 & ~n_21093;
assign n_21095 =  x_300 & ~n_20914;
assign n_21096 =  i_2 &  n_20914;
assign n_21097 = ~n_21095 & ~n_21096;
assign n_21098 =  x_300 & ~n_21097;
assign n_21099 = ~x_300 &  n_21097;
assign n_21100 = ~n_21098 & ~n_21099;
assign n_21101 =  x_299 & ~n_20914;
assign n_21102 =  i_1 &  n_20914;
assign n_21103 = ~n_21101 & ~n_21102;
assign n_21104 =  x_299 & ~n_21103;
assign n_21105 = ~x_299 &  n_21103;
assign n_21106 = ~n_21104 & ~n_21105;
assign n_21107 =  n_3858 &  n_4251;
assign n_21108 =  x_298 & ~n_21107;
assign n_21109 =  i_32 &  n_21107;
assign n_21110 = ~n_21108 & ~n_21109;
assign n_21111 =  x_298 & ~n_21110;
assign n_21112 = ~x_298 &  n_21110;
assign n_21113 = ~n_21111 & ~n_21112;
assign n_21114 =  x_297 & ~n_21107;
assign n_21115 =  i_31 &  n_21107;
assign n_21116 = ~n_21114 & ~n_21115;
assign n_21117 =  x_297 & ~n_21116;
assign n_21118 = ~x_297 &  n_21116;
assign n_21119 = ~n_21117 & ~n_21118;
assign n_21120 =  x_296 & ~n_21107;
assign n_21121 =  i_30 &  n_21107;
assign n_21122 = ~n_21120 & ~n_21121;
assign n_21123 =  x_296 & ~n_21122;
assign n_21124 = ~x_296 &  n_21122;
assign n_21125 = ~n_21123 & ~n_21124;
assign n_21126 =  x_295 & ~n_21107;
assign n_21127 =  i_29 &  n_21107;
assign n_21128 = ~n_21126 & ~n_21127;
assign n_21129 =  x_295 & ~n_21128;
assign n_21130 = ~x_295 &  n_21128;
assign n_21131 = ~n_21129 & ~n_21130;
assign n_21132 =  x_294 & ~n_21107;
assign n_21133 =  i_28 &  n_21107;
assign n_21134 = ~n_21132 & ~n_21133;
assign n_21135 =  x_294 & ~n_21134;
assign n_21136 = ~x_294 &  n_21134;
assign n_21137 = ~n_21135 & ~n_21136;
assign n_21138 =  x_293 & ~n_21107;
assign n_21139 =  i_27 &  n_21107;
assign n_21140 = ~n_21138 & ~n_21139;
assign n_21141 =  x_293 & ~n_21140;
assign n_21142 = ~x_293 &  n_21140;
assign n_21143 = ~n_21141 & ~n_21142;
assign n_21144 =  x_292 & ~n_21107;
assign n_21145 =  i_26 &  n_21107;
assign n_21146 = ~n_21144 & ~n_21145;
assign n_21147 =  x_292 & ~n_21146;
assign n_21148 = ~x_292 &  n_21146;
assign n_21149 = ~n_21147 & ~n_21148;
assign n_21150 =  x_291 & ~n_21107;
assign n_21151 =  i_25 &  n_21107;
assign n_21152 = ~n_21150 & ~n_21151;
assign n_21153 =  x_291 & ~n_21152;
assign n_21154 = ~x_291 &  n_21152;
assign n_21155 = ~n_21153 & ~n_21154;
assign n_21156 =  x_290 & ~n_21107;
assign n_21157 =  i_24 &  n_21107;
assign n_21158 = ~n_21156 & ~n_21157;
assign n_21159 =  x_290 & ~n_21158;
assign n_21160 = ~x_290 &  n_21158;
assign n_21161 = ~n_21159 & ~n_21160;
assign n_21162 =  x_289 & ~n_21107;
assign n_21163 =  i_23 &  n_21107;
assign n_21164 = ~n_21162 & ~n_21163;
assign n_21165 =  x_289 & ~n_21164;
assign n_21166 = ~x_289 &  n_21164;
assign n_21167 = ~n_21165 & ~n_21166;
assign n_21168 =  x_288 & ~n_21107;
assign n_21169 =  i_22 &  n_21107;
assign n_21170 = ~n_21168 & ~n_21169;
assign n_21171 =  x_288 & ~n_21170;
assign n_21172 = ~x_288 &  n_21170;
assign n_21173 = ~n_21171 & ~n_21172;
assign n_21174 =  x_287 & ~n_21107;
assign n_21175 =  i_21 &  n_21107;
assign n_21176 = ~n_21174 & ~n_21175;
assign n_21177 =  x_287 & ~n_21176;
assign n_21178 = ~x_287 &  n_21176;
assign n_21179 = ~n_21177 & ~n_21178;
assign n_21180 =  x_286 & ~n_21107;
assign n_21181 =  i_20 &  n_21107;
assign n_21182 = ~n_21180 & ~n_21181;
assign n_21183 =  x_286 & ~n_21182;
assign n_21184 = ~x_286 &  n_21182;
assign n_21185 = ~n_21183 & ~n_21184;
assign n_21186 =  x_285 & ~n_21107;
assign n_21187 =  i_19 &  n_21107;
assign n_21188 = ~n_21186 & ~n_21187;
assign n_21189 =  x_285 & ~n_21188;
assign n_21190 = ~x_285 &  n_21188;
assign n_21191 = ~n_21189 & ~n_21190;
assign n_21192 =  x_284 & ~n_21107;
assign n_21193 =  i_18 &  n_21107;
assign n_21194 = ~n_21192 & ~n_21193;
assign n_21195 =  x_284 & ~n_21194;
assign n_21196 = ~x_284 &  n_21194;
assign n_21197 = ~n_21195 & ~n_21196;
assign n_21198 =  x_283 & ~n_21107;
assign n_21199 =  i_17 &  n_21107;
assign n_21200 = ~n_21198 & ~n_21199;
assign n_21201 =  x_283 & ~n_21200;
assign n_21202 = ~x_283 &  n_21200;
assign n_21203 = ~n_21201 & ~n_21202;
assign n_21204 =  x_282 & ~n_21107;
assign n_21205 =  i_16 &  n_21107;
assign n_21206 = ~n_21204 & ~n_21205;
assign n_21207 =  x_282 & ~n_21206;
assign n_21208 = ~x_282 &  n_21206;
assign n_21209 = ~n_21207 & ~n_21208;
assign n_21210 =  x_281 & ~n_21107;
assign n_21211 =  i_15 &  n_21107;
assign n_21212 = ~n_21210 & ~n_21211;
assign n_21213 =  x_281 & ~n_21212;
assign n_21214 = ~x_281 &  n_21212;
assign n_21215 = ~n_21213 & ~n_21214;
assign n_21216 =  x_280 & ~n_21107;
assign n_21217 =  i_14 &  n_21107;
assign n_21218 = ~n_21216 & ~n_21217;
assign n_21219 =  x_280 & ~n_21218;
assign n_21220 = ~x_280 &  n_21218;
assign n_21221 = ~n_21219 & ~n_21220;
assign n_21222 =  x_279 & ~n_21107;
assign n_21223 =  i_13 &  n_21107;
assign n_21224 = ~n_21222 & ~n_21223;
assign n_21225 =  x_279 & ~n_21224;
assign n_21226 = ~x_279 &  n_21224;
assign n_21227 = ~n_21225 & ~n_21226;
assign n_21228 =  x_278 & ~n_21107;
assign n_21229 =  i_12 &  n_21107;
assign n_21230 = ~n_21228 & ~n_21229;
assign n_21231 =  x_278 & ~n_21230;
assign n_21232 = ~x_278 &  n_21230;
assign n_21233 = ~n_21231 & ~n_21232;
assign n_21234 =  x_277 & ~n_21107;
assign n_21235 =  i_11 &  n_21107;
assign n_21236 = ~n_21234 & ~n_21235;
assign n_21237 =  x_277 & ~n_21236;
assign n_21238 = ~x_277 &  n_21236;
assign n_21239 = ~n_21237 & ~n_21238;
assign n_21240 =  x_276 & ~n_21107;
assign n_21241 =  i_10 &  n_21107;
assign n_21242 = ~n_21240 & ~n_21241;
assign n_21243 =  x_276 & ~n_21242;
assign n_21244 = ~x_276 &  n_21242;
assign n_21245 = ~n_21243 & ~n_21244;
assign n_21246 =  x_275 & ~n_21107;
assign n_21247 =  i_9 &  n_21107;
assign n_21248 = ~n_21246 & ~n_21247;
assign n_21249 =  x_275 & ~n_21248;
assign n_21250 = ~x_275 &  n_21248;
assign n_21251 = ~n_21249 & ~n_21250;
assign n_21252 =  x_274 & ~n_21107;
assign n_21253 =  i_8 &  n_21107;
assign n_21254 = ~n_21252 & ~n_21253;
assign n_21255 =  x_274 & ~n_21254;
assign n_21256 = ~x_274 &  n_21254;
assign n_21257 = ~n_21255 & ~n_21256;
assign n_21258 =  x_273 & ~n_21107;
assign n_21259 =  i_7 &  n_21107;
assign n_21260 = ~n_21258 & ~n_21259;
assign n_21261 =  x_273 & ~n_21260;
assign n_21262 = ~x_273 &  n_21260;
assign n_21263 = ~n_21261 & ~n_21262;
assign n_21264 =  x_272 & ~n_21107;
assign n_21265 =  i_6 &  n_21107;
assign n_21266 = ~n_21264 & ~n_21265;
assign n_21267 =  x_272 & ~n_21266;
assign n_21268 = ~x_272 &  n_21266;
assign n_21269 = ~n_21267 & ~n_21268;
assign n_21270 =  x_271 & ~n_21107;
assign n_21271 =  i_5 &  n_21107;
assign n_21272 = ~n_21270 & ~n_21271;
assign n_21273 =  x_271 & ~n_21272;
assign n_21274 = ~x_271 &  n_21272;
assign n_21275 = ~n_21273 & ~n_21274;
assign n_21276 =  x_270 & ~n_21107;
assign n_21277 =  i_4 &  n_21107;
assign n_21278 = ~n_21276 & ~n_21277;
assign n_21279 =  x_270 & ~n_21278;
assign n_21280 = ~x_270 &  n_21278;
assign n_21281 = ~n_21279 & ~n_21280;
assign n_21282 =  x_269 & ~n_21107;
assign n_21283 =  i_3 &  n_21107;
assign n_21284 = ~n_21282 & ~n_21283;
assign n_21285 =  x_269 & ~n_21284;
assign n_21286 = ~x_269 &  n_21284;
assign n_21287 = ~n_21285 & ~n_21286;
assign n_21288 =  x_268 & ~n_21107;
assign n_21289 =  i_2 &  n_21107;
assign n_21290 = ~n_21288 & ~n_21289;
assign n_21291 =  x_268 & ~n_21290;
assign n_21292 = ~x_268 &  n_21290;
assign n_21293 = ~n_21291 & ~n_21292;
assign n_21294 =  x_267 & ~n_21107;
assign n_21295 =  i_1 &  n_21107;
assign n_21296 = ~n_21294 & ~n_21295;
assign n_21297 =  x_267 & ~n_21296;
assign n_21298 = ~x_267 &  n_21296;
assign n_21299 = ~n_21297 & ~n_21298;
assign n_21300 =  n_980 &  n_4057;
assign n_21301 =  x_266 & ~n_21300;
assign n_21302 =  i_32 &  n_21300;
assign n_21303 = ~n_21301 & ~n_21302;
assign n_21304 =  x_266 & ~n_21303;
assign n_21305 = ~x_266 &  n_21303;
assign n_21306 = ~n_21304 & ~n_21305;
assign n_21307 =  x_265 & ~n_21300;
assign n_21308 =  i_31 &  n_21300;
assign n_21309 = ~n_21307 & ~n_21308;
assign n_21310 =  x_265 & ~n_21309;
assign n_21311 = ~x_265 &  n_21309;
assign n_21312 = ~n_21310 & ~n_21311;
assign n_21313 =  x_264 & ~n_21300;
assign n_21314 =  i_30 &  n_21300;
assign n_21315 = ~n_21313 & ~n_21314;
assign n_21316 =  x_264 & ~n_21315;
assign n_21317 = ~x_264 &  n_21315;
assign n_21318 = ~n_21316 & ~n_21317;
assign n_21319 =  x_263 & ~n_21300;
assign n_21320 =  i_29 &  n_21300;
assign n_21321 = ~n_21319 & ~n_21320;
assign n_21322 =  x_263 & ~n_21321;
assign n_21323 = ~x_263 &  n_21321;
assign n_21324 = ~n_21322 & ~n_21323;
assign n_21325 =  x_262 & ~n_21300;
assign n_21326 =  i_28 &  n_21300;
assign n_21327 = ~n_21325 & ~n_21326;
assign n_21328 =  x_262 & ~n_21327;
assign n_21329 = ~x_262 &  n_21327;
assign n_21330 = ~n_21328 & ~n_21329;
assign n_21331 =  x_261 & ~n_21300;
assign n_21332 =  i_27 &  n_21300;
assign n_21333 = ~n_21331 & ~n_21332;
assign n_21334 =  x_261 & ~n_21333;
assign n_21335 = ~x_261 &  n_21333;
assign n_21336 = ~n_21334 & ~n_21335;
assign n_21337 =  x_260 & ~n_21300;
assign n_21338 =  i_26 &  n_21300;
assign n_21339 = ~n_21337 & ~n_21338;
assign n_21340 =  x_260 & ~n_21339;
assign n_21341 = ~x_260 &  n_21339;
assign n_21342 = ~n_21340 & ~n_21341;
assign n_21343 =  x_259 & ~n_21300;
assign n_21344 =  i_25 &  n_21300;
assign n_21345 = ~n_21343 & ~n_21344;
assign n_21346 =  x_259 & ~n_21345;
assign n_21347 = ~x_259 &  n_21345;
assign n_21348 = ~n_21346 & ~n_21347;
assign n_21349 =  x_258 & ~n_21300;
assign n_21350 =  i_24 &  n_21300;
assign n_21351 = ~n_21349 & ~n_21350;
assign n_21352 =  x_258 & ~n_21351;
assign n_21353 = ~x_258 &  n_21351;
assign n_21354 = ~n_21352 & ~n_21353;
assign n_21355 =  x_257 & ~n_21300;
assign n_21356 =  i_23 &  n_21300;
assign n_21357 = ~n_21355 & ~n_21356;
assign n_21358 =  x_257 & ~n_21357;
assign n_21359 = ~x_257 &  n_21357;
assign n_21360 = ~n_21358 & ~n_21359;
assign n_21361 =  x_256 & ~n_21300;
assign n_21362 =  i_22 &  n_21300;
assign n_21363 = ~n_21361 & ~n_21362;
assign n_21364 =  x_256 & ~n_21363;
assign n_21365 = ~x_256 &  n_21363;
assign n_21366 = ~n_21364 & ~n_21365;
assign n_21367 =  x_255 & ~n_21300;
assign n_21368 =  i_21 &  n_21300;
assign n_21369 = ~n_21367 & ~n_21368;
assign n_21370 =  x_255 & ~n_21369;
assign n_21371 = ~x_255 &  n_21369;
assign n_21372 = ~n_21370 & ~n_21371;
assign n_21373 =  x_254 & ~n_21300;
assign n_21374 =  i_20 &  n_21300;
assign n_21375 = ~n_21373 & ~n_21374;
assign n_21376 =  x_254 & ~n_21375;
assign n_21377 = ~x_254 &  n_21375;
assign n_21378 = ~n_21376 & ~n_21377;
assign n_21379 =  x_253 & ~n_21300;
assign n_21380 =  i_19 &  n_21300;
assign n_21381 = ~n_21379 & ~n_21380;
assign n_21382 =  x_253 & ~n_21381;
assign n_21383 = ~x_253 &  n_21381;
assign n_21384 = ~n_21382 & ~n_21383;
assign n_21385 =  x_252 & ~n_21300;
assign n_21386 =  i_18 &  n_21300;
assign n_21387 = ~n_21385 & ~n_21386;
assign n_21388 =  x_252 & ~n_21387;
assign n_21389 = ~x_252 &  n_21387;
assign n_21390 = ~n_21388 & ~n_21389;
assign n_21391 =  x_251 & ~n_21300;
assign n_21392 =  i_17 &  n_21300;
assign n_21393 = ~n_21391 & ~n_21392;
assign n_21394 =  x_251 & ~n_21393;
assign n_21395 = ~x_251 &  n_21393;
assign n_21396 = ~n_21394 & ~n_21395;
assign n_21397 =  x_250 & ~n_21300;
assign n_21398 =  i_16 &  n_21300;
assign n_21399 = ~n_21397 & ~n_21398;
assign n_21400 =  x_250 & ~n_21399;
assign n_21401 = ~x_250 &  n_21399;
assign n_21402 = ~n_21400 & ~n_21401;
assign n_21403 =  x_249 & ~n_21300;
assign n_21404 =  i_15 &  n_21300;
assign n_21405 = ~n_21403 & ~n_21404;
assign n_21406 =  x_249 & ~n_21405;
assign n_21407 = ~x_249 &  n_21405;
assign n_21408 = ~n_21406 & ~n_21407;
assign n_21409 =  x_248 & ~n_21300;
assign n_21410 =  i_14 &  n_21300;
assign n_21411 = ~n_21409 & ~n_21410;
assign n_21412 =  x_248 & ~n_21411;
assign n_21413 = ~x_248 &  n_21411;
assign n_21414 = ~n_21412 & ~n_21413;
assign n_21415 =  x_247 & ~n_21300;
assign n_21416 =  i_13 &  n_21300;
assign n_21417 = ~n_21415 & ~n_21416;
assign n_21418 =  x_247 & ~n_21417;
assign n_21419 = ~x_247 &  n_21417;
assign n_21420 = ~n_21418 & ~n_21419;
assign n_21421 =  x_246 & ~n_21300;
assign n_21422 =  i_12 &  n_21300;
assign n_21423 = ~n_21421 & ~n_21422;
assign n_21424 =  x_246 & ~n_21423;
assign n_21425 = ~x_246 &  n_21423;
assign n_21426 = ~n_21424 & ~n_21425;
assign n_21427 =  x_245 & ~n_21300;
assign n_21428 =  i_11 &  n_21300;
assign n_21429 = ~n_21427 & ~n_21428;
assign n_21430 =  x_245 & ~n_21429;
assign n_21431 = ~x_245 &  n_21429;
assign n_21432 = ~n_21430 & ~n_21431;
assign n_21433 =  x_244 & ~n_21300;
assign n_21434 =  i_10 &  n_21300;
assign n_21435 = ~n_21433 & ~n_21434;
assign n_21436 =  x_244 & ~n_21435;
assign n_21437 = ~x_244 &  n_21435;
assign n_21438 = ~n_21436 & ~n_21437;
assign n_21439 =  x_243 & ~n_21300;
assign n_21440 =  i_9 &  n_21300;
assign n_21441 = ~n_21439 & ~n_21440;
assign n_21442 =  x_243 & ~n_21441;
assign n_21443 = ~x_243 &  n_21441;
assign n_21444 = ~n_21442 & ~n_21443;
assign n_21445 =  x_242 & ~n_21300;
assign n_21446 =  i_8 &  n_21300;
assign n_21447 = ~n_21445 & ~n_21446;
assign n_21448 =  x_242 & ~n_21447;
assign n_21449 = ~x_242 &  n_21447;
assign n_21450 = ~n_21448 & ~n_21449;
assign n_21451 =  x_241 & ~n_21300;
assign n_21452 =  i_7 &  n_21300;
assign n_21453 = ~n_21451 & ~n_21452;
assign n_21454 =  x_241 & ~n_21453;
assign n_21455 = ~x_241 &  n_21453;
assign n_21456 = ~n_21454 & ~n_21455;
assign n_21457 =  x_240 & ~n_21300;
assign n_21458 =  i_6 &  n_21300;
assign n_21459 = ~n_21457 & ~n_21458;
assign n_21460 =  x_240 & ~n_21459;
assign n_21461 = ~x_240 &  n_21459;
assign n_21462 = ~n_21460 & ~n_21461;
assign n_21463 =  x_239 & ~n_21300;
assign n_21464 =  i_5 &  n_21300;
assign n_21465 = ~n_21463 & ~n_21464;
assign n_21466 =  x_239 & ~n_21465;
assign n_21467 = ~x_239 &  n_21465;
assign n_21468 = ~n_21466 & ~n_21467;
assign n_21469 =  x_238 & ~n_21300;
assign n_21470 =  i_4 &  n_21300;
assign n_21471 = ~n_21469 & ~n_21470;
assign n_21472 =  x_238 & ~n_21471;
assign n_21473 = ~x_238 &  n_21471;
assign n_21474 = ~n_21472 & ~n_21473;
assign n_21475 =  x_237 & ~n_21300;
assign n_21476 =  i_3 &  n_21300;
assign n_21477 = ~n_21475 & ~n_21476;
assign n_21478 =  x_237 & ~n_21477;
assign n_21479 = ~x_237 &  n_21477;
assign n_21480 = ~n_21478 & ~n_21479;
assign n_21481 =  x_236 & ~n_21300;
assign n_21482 =  i_2 &  n_21300;
assign n_21483 = ~n_21481 & ~n_21482;
assign n_21484 =  x_236 & ~n_21483;
assign n_21485 = ~x_236 &  n_21483;
assign n_21486 = ~n_21484 & ~n_21485;
assign n_21487 =  x_235 & ~n_21300;
assign n_21488 =  i_1 &  n_21300;
assign n_21489 = ~n_21487 & ~n_21488;
assign n_21490 =  x_235 & ~n_21489;
assign n_21491 = ~x_235 &  n_21489;
assign n_21492 = ~n_21490 & ~n_21491;
assign n_21493 =  n_3 &  n_191;
assign n_21494 =  x_234 & ~n_21493;
assign n_21495 =  i_32 &  n_21493;
assign n_21496 = ~n_21494 & ~n_21495;
assign n_21497 =  x_234 & ~n_21496;
assign n_21498 = ~x_234 &  n_21496;
assign n_21499 = ~n_21497 & ~n_21498;
assign n_21500 =  x_233 & ~n_21493;
assign n_21501 =  i_31 &  n_21493;
assign n_21502 = ~n_21500 & ~n_21501;
assign n_21503 =  x_233 & ~n_21502;
assign n_21504 = ~x_233 &  n_21502;
assign n_21505 = ~n_21503 & ~n_21504;
assign n_21506 =  x_232 & ~n_21493;
assign n_21507 =  i_30 &  n_21493;
assign n_21508 = ~n_21506 & ~n_21507;
assign n_21509 =  x_232 & ~n_21508;
assign n_21510 = ~x_232 &  n_21508;
assign n_21511 = ~n_21509 & ~n_21510;
assign n_21512 =  x_231 & ~n_21493;
assign n_21513 =  i_29 &  n_21493;
assign n_21514 = ~n_21512 & ~n_21513;
assign n_21515 =  x_231 & ~n_21514;
assign n_21516 = ~x_231 &  n_21514;
assign n_21517 = ~n_21515 & ~n_21516;
assign n_21518 =  x_230 & ~n_21493;
assign n_21519 =  i_28 &  n_21493;
assign n_21520 = ~n_21518 & ~n_21519;
assign n_21521 =  x_230 & ~n_21520;
assign n_21522 = ~x_230 &  n_21520;
assign n_21523 = ~n_21521 & ~n_21522;
assign n_21524 =  x_229 & ~n_21493;
assign n_21525 =  i_27 &  n_21493;
assign n_21526 = ~n_21524 & ~n_21525;
assign n_21527 =  x_229 & ~n_21526;
assign n_21528 = ~x_229 &  n_21526;
assign n_21529 = ~n_21527 & ~n_21528;
assign n_21530 =  x_228 & ~n_21493;
assign n_21531 =  i_26 &  n_21493;
assign n_21532 = ~n_21530 & ~n_21531;
assign n_21533 =  x_228 & ~n_21532;
assign n_21534 = ~x_228 &  n_21532;
assign n_21535 = ~n_21533 & ~n_21534;
assign n_21536 =  x_227 & ~n_21493;
assign n_21537 =  i_25 &  n_21493;
assign n_21538 = ~n_21536 & ~n_21537;
assign n_21539 =  x_227 & ~n_21538;
assign n_21540 = ~x_227 &  n_21538;
assign n_21541 = ~n_21539 & ~n_21540;
assign n_21542 =  x_226 & ~n_21493;
assign n_21543 =  i_24 &  n_21493;
assign n_21544 = ~n_21542 & ~n_21543;
assign n_21545 =  x_226 & ~n_21544;
assign n_21546 = ~x_226 &  n_21544;
assign n_21547 = ~n_21545 & ~n_21546;
assign n_21548 =  x_225 & ~n_21493;
assign n_21549 =  i_23 &  n_21493;
assign n_21550 = ~n_21548 & ~n_21549;
assign n_21551 =  x_225 & ~n_21550;
assign n_21552 = ~x_225 &  n_21550;
assign n_21553 = ~n_21551 & ~n_21552;
assign n_21554 =  x_224 & ~n_21493;
assign n_21555 =  i_22 &  n_21493;
assign n_21556 = ~n_21554 & ~n_21555;
assign n_21557 =  x_224 & ~n_21556;
assign n_21558 = ~x_224 &  n_21556;
assign n_21559 = ~n_21557 & ~n_21558;
assign n_21560 =  x_223 & ~n_21493;
assign n_21561 =  i_21 &  n_21493;
assign n_21562 = ~n_21560 & ~n_21561;
assign n_21563 =  x_223 & ~n_21562;
assign n_21564 = ~x_223 &  n_21562;
assign n_21565 = ~n_21563 & ~n_21564;
assign n_21566 =  x_222 & ~n_21493;
assign n_21567 =  i_20 &  n_21493;
assign n_21568 = ~n_21566 & ~n_21567;
assign n_21569 =  x_222 & ~n_21568;
assign n_21570 = ~x_222 &  n_21568;
assign n_21571 = ~n_21569 & ~n_21570;
assign n_21572 =  x_221 & ~n_21493;
assign n_21573 =  i_19 &  n_21493;
assign n_21574 = ~n_21572 & ~n_21573;
assign n_21575 =  x_221 & ~n_21574;
assign n_21576 = ~x_221 &  n_21574;
assign n_21577 = ~n_21575 & ~n_21576;
assign n_21578 =  x_220 & ~n_21493;
assign n_21579 =  i_18 &  n_21493;
assign n_21580 = ~n_21578 & ~n_21579;
assign n_21581 =  x_220 & ~n_21580;
assign n_21582 = ~x_220 &  n_21580;
assign n_21583 = ~n_21581 & ~n_21582;
assign n_21584 =  x_219 & ~n_21493;
assign n_21585 =  i_17 &  n_21493;
assign n_21586 = ~n_21584 & ~n_21585;
assign n_21587 =  x_219 & ~n_21586;
assign n_21588 = ~x_219 &  n_21586;
assign n_21589 = ~n_21587 & ~n_21588;
assign n_21590 =  x_218 & ~n_21493;
assign n_21591 =  i_16 &  n_21493;
assign n_21592 = ~n_21590 & ~n_21591;
assign n_21593 =  x_218 & ~n_21592;
assign n_21594 = ~x_218 &  n_21592;
assign n_21595 = ~n_21593 & ~n_21594;
assign n_21596 =  x_217 & ~n_21493;
assign n_21597 =  i_15 &  n_21493;
assign n_21598 = ~n_21596 & ~n_21597;
assign n_21599 =  x_217 & ~n_21598;
assign n_21600 = ~x_217 &  n_21598;
assign n_21601 = ~n_21599 & ~n_21600;
assign n_21602 =  x_216 & ~n_21493;
assign n_21603 =  i_14 &  n_21493;
assign n_21604 = ~n_21602 & ~n_21603;
assign n_21605 =  x_216 & ~n_21604;
assign n_21606 = ~x_216 &  n_21604;
assign n_21607 = ~n_21605 & ~n_21606;
assign n_21608 =  x_215 & ~n_21493;
assign n_21609 =  i_13 &  n_21493;
assign n_21610 = ~n_21608 & ~n_21609;
assign n_21611 =  x_215 & ~n_21610;
assign n_21612 = ~x_215 &  n_21610;
assign n_21613 = ~n_21611 & ~n_21612;
assign n_21614 =  x_214 & ~n_21493;
assign n_21615 =  i_12 &  n_21493;
assign n_21616 = ~n_21614 & ~n_21615;
assign n_21617 =  x_214 & ~n_21616;
assign n_21618 = ~x_214 &  n_21616;
assign n_21619 = ~n_21617 & ~n_21618;
assign n_21620 =  x_213 & ~n_21493;
assign n_21621 =  i_11 &  n_21493;
assign n_21622 = ~n_21620 & ~n_21621;
assign n_21623 =  x_213 & ~n_21622;
assign n_21624 = ~x_213 &  n_21622;
assign n_21625 = ~n_21623 & ~n_21624;
assign n_21626 =  x_212 & ~n_21493;
assign n_21627 =  i_10 &  n_21493;
assign n_21628 = ~n_21626 & ~n_21627;
assign n_21629 =  x_212 & ~n_21628;
assign n_21630 = ~x_212 &  n_21628;
assign n_21631 = ~n_21629 & ~n_21630;
assign n_21632 =  x_211 & ~n_21493;
assign n_21633 =  i_9 &  n_21493;
assign n_21634 = ~n_21632 & ~n_21633;
assign n_21635 =  x_211 & ~n_21634;
assign n_21636 = ~x_211 &  n_21634;
assign n_21637 = ~n_21635 & ~n_21636;
assign n_21638 =  x_210 & ~n_21493;
assign n_21639 =  i_8 &  n_21493;
assign n_21640 = ~n_21638 & ~n_21639;
assign n_21641 =  x_210 & ~n_21640;
assign n_21642 = ~x_210 &  n_21640;
assign n_21643 = ~n_21641 & ~n_21642;
assign n_21644 =  x_209 & ~n_21493;
assign n_21645 =  i_7 &  n_21493;
assign n_21646 = ~n_21644 & ~n_21645;
assign n_21647 =  x_209 & ~n_21646;
assign n_21648 = ~x_209 &  n_21646;
assign n_21649 = ~n_21647 & ~n_21648;
assign n_21650 =  x_208 & ~n_21493;
assign n_21651 =  i_6 &  n_21493;
assign n_21652 = ~n_21650 & ~n_21651;
assign n_21653 =  x_208 & ~n_21652;
assign n_21654 = ~x_208 &  n_21652;
assign n_21655 = ~n_21653 & ~n_21654;
assign n_21656 =  x_207 & ~n_21493;
assign n_21657 =  i_5 &  n_21493;
assign n_21658 = ~n_21656 & ~n_21657;
assign n_21659 =  x_207 & ~n_21658;
assign n_21660 = ~x_207 &  n_21658;
assign n_21661 = ~n_21659 & ~n_21660;
assign n_21662 =  x_206 & ~n_21493;
assign n_21663 =  i_4 &  n_21493;
assign n_21664 = ~n_21662 & ~n_21663;
assign n_21665 =  x_206 & ~n_21664;
assign n_21666 = ~x_206 &  n_21664;
assign n_21667 = ~n_21665 & ~n_21666;
assign n_21668 =  x_205 & ~n_21493;
assign n_21669 =  i_3 &  n_21493;
assign n_21670 = ~n_21668 & ~n_21669;
assign n_21671 =  x_205 & ~n_21670;
assign n_21672 = ~x_205 &  n_21670;
assign n_21673 = ~n_21671 & ~n_21672;
assign n_21674 =  x_204 & ~n_21493;
assign n_21675 =  i_2 &  n_21493;
assign n_21676 = ~n_21674 & ~n_21675;
assign n_21677 =  x_204 & ~n_21676;
assign n_21678 = ~x_204 &  n_21676;
assign n_21679 = ~n_21677 & ~n_21678;
assign n_21680 =  x_203 & ~n_21493;
assign n_21681 =  i_1 &  n_21493;
assign n_21682 = ~n_21680 & ~n_21681;
assign n_21683 =  x_203 & ~n_21682;
assign n_21684 = ~x_203 &  n_21682;
assign n_21685 = ~n_21683 & ~n_21684;
assign n_21686 =  n_4993 &  n_3275;
assign n_21687 =  x_202 & ~n_21686;
assign n_21688 =  i_32 &  n_21686;
assign n_21689 = ~n_21687 & ~n_21688;
assign n_21690 =  x_202 & ~n_21689;
assign n_21691 = ~x_202 &  n_21689;
assign n_21692 = ~n_21690 & ~n_21691;
assign n_21693 =  x_201 & ~n_21686;
assign n_21694 =  i_31 &  n_21686;
assign n_21695 = ~n_21693 & ~n_21694;
assign n_21696 =  x_201 & ~n_21695;
assign n_21697 = ~x_201 &  n_21695;
assign n_21698 = ~n_21696 & ~n_21697;
assign n_21699 =  x_200 & ~n_21686;
assign n_21700 =  i_30 &  n_21686;
assign n_21701 = ~n_21699 & ~n_21700;
assign n_21702 =  x_200 & ~n_21701;
assign n_21703 = ~x_200 &  n_21701;
assign n_21704 = ~n_21702 & ~n_21703;
assign n_21705 =  x_199 & ~n_21686;
assign n_21706 =  i_29 &  n_21686;
assign n_21707 = ~n_21705 & ~n_21706;
assign n_21708 =  x_199 & ~n_21707;
assign n_21709 = ~x_199 &  n_21707;
assign n_21710 = ~n_21708 & ~n_21709;
assign n_21711 =  x_198 & ~n_21686;
assign n_21712 =  i_28 &  n_21686;
assign n_21713 = ~n_21711 & ~n_21712;
assign n_21714 =  x_198 & ~n_21713;
assign n_21715 = ~x_198 &  n_21713;
assign n_21716 = ~n_21714 & ~n_21715;
assign n_21717 =  x_197 & ~n_21686;
assign n_21718 =  i_27 &  n_21686;
assign n_21719 = ~n_21717 & ~n_21718;
assign n_21720 =  x_197 & ~n_21719;
assign n_21721 = ~x_197 &  n_21719;
assign n_21722 = ~n_21720 & ~n_21721;
assign n_21723 =  x_196 & ~n_21686;
assign n_21724 =  i_26 &  n_21686;
assign n_21725 = ~n_21723 & ~n_21724;
assign n_21726 =  x_196 & ~n_21725;
assign n_21727 = ~x_196 &  n_21725;
assign n_21728 = ~n_21726 & ~n_21727;
assign n_21729 =  x_195 & ~n_21686;
assign n_21730 =  i_25 &  n_21686;
assign n_21731 = ~n_21729 & ~n_21730;
assign n_21732 =  x_195 & ~n_21731;
assign n_21733 = ~x_195 &  n_21731;
assign n_21734 = ~n_21732 & ~n_21733;
assign n_21735 =  x_194 & ~n_21686;
assign n_21736 =  i_24 &  n_21686;
assign n_21737 = ~n_21735 & ~n_21736;
assign n_21738 =  x_194 & ~n_21737;
assign n_21739 = ~x_194 &  n_21737;
assign n_21740 = ~n_21738 & ~n_21739;
assign n_21741 =  x_193 & ~n_21686;
assign n_21742 =  i_23 &  n_21686;
assign n_21743 = ~n_21741 & ~n_21742;
assign n_21744 =  x_193 & ~n_21743;
assign n_21745 = ~x_193 &  n_21743;
assign n_21746 = ~n_21744 & ~n_21745;
assign n_21747 =  x_192 & ~n_21686;
assign n_21748 =  i_22 &  n_21686;
assign n_21749 = ~n_21747 & ~n_21748;
assign n_21750 =  x_192 & ~n_21749;
assign n_21751 = ~x_192 &  n_21749;
assign n_21752 = ~n_21750 & ~n_21751;
assign n_21753 =  x_191 & ~n_21686;
assign n_21754 =  i_21 &  n_21686;
assign n_21755 = ~n_21753 & ~n_21754;
assign n_21756 =  x_191 & ~n_21755;
assign n_21757 = ~x_191 &  n_21755;
assign n_21758 = ~n_21756 & ~n_21757;
assign n_21759 =  x_190 & ~n_21686;
assign n_21760 =  i_20 &  n_21686;
assign n_21761 = ~n_21759 & ~n_21760;
assign n_21762 =  x_190 & ~n_21761;
assign n_21763 = ~x_190 &  n_21761;
assign n_21764 = ~n_21762 & ~n_21763;
assign n_21765 =  x_189 & ~n_21686;
assign n_21766 =  i_19 &  n_21686;
assign n_21767 = ~n_21765 & ~n_21766;
assign n_21768 =  x_189 & ~n_21767;
assign n_21769 = ~x_189 &  n_21767;
assign n_21770 = ~n_21768 & ~n_21769;
assign n_21771 =  x_188 & ~n_21686;
assign n_21772 =  i_18 &  n_21686;
assign n_21773 = ~n_21771 & ~n_21772;
assign n_21774 =  x_188 & ~n_21773;
assign n_21775 = ~x_188 &  n_21773;
assign n_21776 = ~n_21774 & ~n_21775;
assign n_21777 =  x_187 & ~n_21686;
assign n_21778 =  i_17 &  n_21686;
assign n_21779 = ~n_21777 & ~n_21778;
assign n_21780 =  x_187 & ~n_21779;
assign n_21781 = ~x_187 &  n_21779;
assign n_21782 = ~n_21780 & ~n_21781;
assign n_21783 =  x_186 & ~n_21686;
assign n_21784 =  i_16 &  n_21686;
assign n_21785 = ~n_21783 & ~n_21784;
assign n_21786 =  x_186 & ~n_21785;
assign n_21787 = ~x_186 &  n_21785;
assign n_21788 = ~n_21786 & ~n_21787;
assign n_21789 =  x_185 & ~n_21686;
assign n_21790 =  i_15 &  n_21686;
assign n_21791 = ~n_21789 & ~n_21790;
assign n_21792 =  x_185 & ~n_21791;
assign n_21793 = ~x_185 &  n_21791;
assign n_21794 = ~n_21792 & ~n_21793;
assign n_21795 =  x_184 & ~n_21686;
assign n_21796 =  i_14 &  n_21686;
assign n_21797 = ~n_21795 & ~n_21796;
assign n_21798 =  x_184 & ~n_21797;
assign n_21799 = ~x_184 &  n_21797;
assign n_21800 = ~n_21798 & ~n_21799;
assign n_21801 =  x_183 & ~n_21686;
assign n_21802 =  i_13 &  n_21686;
assign n_21803 = ~n_21801 & ~n_21802;
assign n_21804 =  x_183 & ~n_21803;
assign n_21805 = ~x_183 &  n_21803;
assign n_21806 = ~n_21804 & ~n_21805;
assign n_21807 =  x_182 & ~n_21686;
assign n_21808 =  i_12 &  n_21686;
assign n_21809 = ~n_21807 & ~n_21808;
assign n_21810 =  x_182 & ~n_21809;
assign n_21811 = ~x_182 &  n_21809;
assign n_21812 = ~n_21810 & ~n_21811;
assign n_21813 =  x_181 & ~n_21686;
assign n_21814 =  i_11 &  n_21686;
assign n_21815 = ~n_21813 & ~n_21814;
assign n_21816 =  x_181 & ~n_21815;
assign n_21817 = ~x_181 &  n_21815;
assign n_21818 = ~n_21816 & ~n_21817;
assign n_21819 =  x_180 & ~n_21686;
assign n_21820 =  i_10 &  n_21686;
assign n_21821 = ~n_21819 & ~n_21820;
assign n_21822 =  x_180 & ~n_21821;
assign n_21823 = ~x_180 &  n_21821;
assign n_21824 = ~n_21822 & ~n_21823;
assign n_21825 =  x_179 & ~n_21686;
assign n_21826 =  i_9 &  n_21686;
assign n_21827 = ~n_21825 & ~n_21826;
assign n_21828 =  x_179 & ~n_21827;
assign n_21829 = ~x_179 &  n_21827;
assign n_21830 = ~n_21828 & ~n_21829;
assign n_21831 =  x_178 & ~n_21686;
assign n_21832 =  i_8 &  n_21686;
assign n_21833 = ~n_21831 & ~n_21832;
assign n_21834 =  x_178 & ~n_21833;
assign n_21835 = ~x_178 &  n_21833;
assign n_21836 = ~n_21834 & ~n_21835;
assign n_21837 =  x_177 & ~n_21686;
assign n_21838 =  i_7 &  n_21686;
assign n_21839 = ~n_21837 & ~n_21838;
assign n_21840 =  x_177 & ~n_21839;
assign n_21841 = ~x_177 &  n_21839;
assign n_21842 = ~n_21840 & ~n_21841;
assign n_21843 =  x_176 & ~n_21686;
assign n_21844 =  i_6 &  n_21686;
assign n_21845 = ~n_21843 & ~n_21844;
assign n_21846 =  x_176 & ~n_21845;
assign n_21847 = ~x_176 &  n_21845;
assign n_21848 = ~n_21846 & ~n_21847;
assign n_21849 =  x_175 & ~n_21686;
assign n_21850 =  i_5 &  n_21686;
assign n_21851 = ~n_21849 & ~n_21850;
assign n_21852 =  x_175 & ~n_21851;
assign n_21853 = ~x_175 &  n_21851;
assign n_21854 = ~n_21852 & ~n_21853;
assign n_21855 =  x_174 & ~n_21686;
assign n_21856 =  i_4 &  n_21686;
assign n_21857 = ~n_21855 & ~n_21856;
assign n_21858 =  x_174 & ~n_21857;
assign n_21859 = ~x_174 &  n_21857;
assign n_21860 = ~n_21858 & ~n_21859;
assign n_21861 =  x_173 & ~n_21686;
assign n_21862 =  i_3 &  n_21686;
assign n_21863 = ~n_21861 & ~n_21862;
assign n_21864 =  x_173 & ~n_21863;
assign n_21865 = ~x_173 &  n_21863;
assign n_21866 = ~n_21864 & ~n_21865;
assign n_21867 =  x_172 & ~n_21686;
assign n_21868 =  i_2 &  n_21686;
assign n_21869 = ~n_21867 & ~n_21868;
assign n_21870 =  x_172 & ~n_21869;
assign n_21871 = ~x_172 &  n_21869;
assign n_21872 = ~n_21870 & ~n_21871;
assign n_21873 =  x_171 & ~n_21686;
assign n_21874 =  i_1 &  n_21686;
assign n_21875 = ~n_21873 & ~n_21874;
assign n_21876 =  x_171 & ~n_21875;
assign n_21877 = ~x_171 &  n_21875;
assign n_21878 = ~n_21876 & ~n_21877;
assign n_21879 =  n_1709 &  n_6533;
assign n_21880 =  x_170 & ~n_21879;
assign n_21881 =  i_32 &  n_21879;
assign n_21882 = ~n_21880 & ~n_21881;
assign n_21883 =  x_170 & ~n_21882;
assign n_21884 = ~x_170 &  n_21882;
assign n_21885 = ~n_21883 & ~n_21884;
assign n_21886 =  x_169 & ~n_21879;
assign n_21887 =  i_31 &  n_21879;
assign n_21888 = ~n_21886 & ~n_21887;
assign n_21889 =  x_169 & ~n_21888;
assign n_21890 = ~x_169 &  n_21888;
assign n_21891 = ~n_21889 & ~n_21890;
assign n_21892 =  x_168 & ~n_21879;
assign n_21893 =  i_30 &  n_21879;
assign n_21894 = ~n_21892 & ~n_21893;
assign n_21895 =  x_168 & ~n_21894;
assign n_21896 = ~x_168 &  n_21894;
assign n_21897 = ~n_21895 & ~n_21896;
assign n_21898 =  x_167 & ~n_21879;
assign n_21899 =  i_29 &  n_21879;
assign n_21900 = ~n_21898 & ~n_21899;
assign n_21901 =  x_167 & ~n_21900;
assign n_21902 = ~x_167 &  n_21900;
assign n_21903 = ~n_21901 & ~n_21902;
assign n_21904 =  x_166 & ~n_21879;
assign n_21905 =  i_28 &  n_21879;
assign n_21906 = ~n_21904 & ~n_21905;
assign n_21907 =  x_166 & ~n_21906;
assign n_21908 = ~x_166 &  n_21906;
assign n_21909 = ~n_21907 & ~n_21908;
assign n_21910 =  x_165 & ~n_21879;
assign n_21911 =  i_27 &  n_21879;
assign n_21912 = ~n_21910 & ~n_21911;
assign n_21913 =  x_165 & ~n_21912;
assign n_21914 = ~x_165 &  n_21912;
assign n_21915 = ~n_21913 & ~n_21914;
assign n_21916 =  x_164 & ~n_21879;
assign n_21917 =  i_26 &  n_21879;
assign n_21918 = ~n_21916 & ~n_21917;
assign n_21919 =  x_164 & ~n_21918;
assign n_21920 = ~x_164 &  n_21918;
assign n_21921 = ~n_21919 & ~n_21920;
assign n_21922 =  x_163 & ~n_21879;
assign n_21923 =  i_25 &  n_21879;
assign n_21924 = ~n_21922 & ~n_21923;
assign n_21925 =  x_163 & ~n_21924;
assign n_21926 = ~x_163 &  n_21924;
assign n_21927 = ~n_21925 & ~n_21926;
assign n_21928 =  x_162 & ~n_21879;
assign n_21929 =  i_24 &  n_21879;
assign n_21930 = ~n_21928 & ~n_21929;
assign n_21931 =  x_162 & ~n_21930;
assign n_21932 = ~x_162 &  n_21930;
assign n_21933 = ~n_21931 & ~n_21932;
assign n_21934 =  x_161 & ~n_21879;
assign n_21935 =  i_23 &  n_21879;
assign n_21936 = ~n_21934 & ~n_21935;
assign n_21937 =  x_161 & ~n_21936;
assign n_21938 = ~x_161 &  n_21936;
assign n_21939 = ~n_21937 & ~n_21938;
assign n_21940 =  x_160 & ~n_21879;
assign n_21941 =  i_22 &  n_21879;
assign n_21942 = ~n_21940 & ~n_21941;
assign n_21943 =  x_160 & ~n_21942;
assign n_21944 = ~x_160 &  n_21942;
assign n_21945 = ~n_21943 & ~n_21944;
assign n_21946 =  x_159 & ~n_21879;
assign n_21947 =  i_21 &  n_21879;
assign n_21948 = ~n_21946 & ~n_21947;
assign n_21949 =  x_159 & ~n_21948;
assign n_21950 = ~x_159 &  n_21948;
assign n_21951 = ~n_21949 & ~n_21950;
assign n_21952 =  x_158 & ~n_21879;
assign n_21953 =  i_20 &  n_21879;
assign n_21954 = ~n_21952 & ~n_21953;
assign n_21955 =  x_158 & ~n_21954;
assign n_21956 = ~x_158 &  n_21954;
assign n_21957 = ~n_21955 & ~n_21956;
assign n_21958 =  x_157 & ~n_21879;
assign n_21959 =  i_19 &  n_21879;
assign n_21960 = ~n_21958 & ~n_21959;
assign n_21961 =  x_157 & ~n_21960;
assign n_21962 = ~x_157 &  n_21960;
assign n_21963 = ~n_21961 & ~n_21962;
assign n_21964 =  x_156 & ~n_21879;
assign n_21965 =  i_18 &  n_21879;
assign n_21966 = ~n_21964 & ~n_21965;
assign n_21967 =  x_156 & ~n_21966;
assign n_21968 = ~x_156 &  n_21966;
assign n_21969 = ~n_21967 & ~n_21968;
assign n_21970 =  x_155 & ~n_21879;
assign n_21971 =  i_17 &  n_21879;
assign n_21972 = ~n_21970 & ~n_21971;
assign n_21973 =  x_155 & ~n_21972;
assign n_21974 = ~x_155 &  n_21972;
assign n_21975 = ~n_21973 & ~n_21974;
assign n_21976 =  x_154 & ~n_21879;
assign n_21977 =  i_16 &  n_21879;
assign n_21978 = ~n_21976 & ~n_21977;
assign n_21979 =  x_154 & ~n_21978;
assign n_21980 = ~x_154 &  n_21978;
assign n_21981 = ~n_21979 & ~n_21980;
assign n_21982 =  x_153 & ~n_21879;
assign n_21983 =  i_15 &  n_21879;
assign n_21984 = ~n_21982 & ~n_21983;
assign n_21985 =  x_153 & ~n_21984;
assign n_21986 = ~x_153 &  n_21984;
assign n_21987 = ~n_21985 & ~n_21986;
assign n_21988 =  x_152 & ~n_21879;
assign n_21989 =  i_14 &  n_21879;
assign n_21990 = ~n_21988 & ~n_21989;
assign n_21991 =  x_152 & ~n_21990;
assign n_21992 = ~x_152 &  n_21990;
assign n_21993 = ~n_21991 & ~n_21992;
assign n_21994 =  x_151 & ~n_21879;
assign n_21995 =  i_13 &  n_21879;
assign n_21996 = ~n_21994 & ~n_21995;
assign n_21997 =  x_151 & ~n_21996;
assign n_21998 = ~x_151 &  n_21996;
assign n_21999 = ~n_21997 & ~n_21998;
assign n_22000 =  x_150 & ~n_21879;
assign n_22001 =  i_12 &  n_21879;
assign n_22002 = ~n_22000 & ~n_22001;
assign n_22003 =  x_150 & ~n_22002;
assign n_22004 = ~x_150 &  n_22002;
assign n_22005 = ~n_22003 & ~n_22004;
assign n_22006 =  x_149 & ~n_21879;
assign n_22007 =  i_11 &  n_21879;
assign n_22008 = ~n_22006 & ~n_22007;
assign n_22009 =  x_149 & ~n_22008;
assign n_22010 = ~x_149 &  n_22008;
assign n_22011 = ~n_22009 & ~n_22010;
assign n_22012 =  x_148 & ~n_21879;
assign n_22013 =  i_10 &  n_21879;
assign n_22014 = ~n_22012 & ~n_22013;
assign n_22015 =  x_148 & ~n_22014;
assign n_22016 = ~x_148 &  n_22014;
assign n_22017 = ~n_22015 & ~n_22016;
assign n_22018 =  x_147 & ~n_21879;
assign n_22019 =  i_9 &  n_21879;
assign n_22020 = ~n_22018 & ~n_22019;
assign n_22021 =  x_147 & ~n_22020;
assign n_22022 = ~x_147 &  n_22020;
assign n_22023 = ~n_22021 & ~n_22022;
assign n_22024 =  x_146 & ~n_21879;
assign n_22025 =  i_8 &  n_21879;
assign n_22026 = ~n_22024 & ~n_22025;
assign n_22027 =  x_146 & ~n_22026;
assign n_22028 = ~x_146 &  n_22026;
assign n_22029 = ~n_22027 & ~n_22028;
assign n_22030 =  x_145 & ~n_21879;
assign n_22031 =  i_7 &  n_21879;
assign n_22032 = ~n_22030 & ~n_22031;
assign n_22033 =  x_145 & ~n_22032;
assign n_22034 = ~x_145 &  n_22032;
assign n_22035 = ~n_22033 & ~n_22034;
assign n_22036 =  x_144 & ~n_21879;
assign n_22037 =  i_6 &  n_21879;
assign n_22038 = ~n_22036 & ~n_22037;
assign n_22039 =  x_144 & ~n_22038;
assign n_22040 = ~x_144 &  n_22038;
assign n_22041 = ~n_22039 & ~n_22040;
assign n_22042 =  x_143 & ~n_21879;
assign n_22043 =  i_5 &  n_21879;
assign n_22044 = ~n_22042 & ~n_22043;
assign n_22045 =  x_143 & ~n_22044;
assign n_22046 = ~x_143 &  n_22044;
assign n_22047 = ~n_22045 & ~n_22046;
assign n_22048 =  x_142 & ~n_21879;
assign n_22049 =  i_4 &  n_21879;
assign n_22050 = ~n_22048 & ~n_22049;
assign n_22051 =  x_142 & ~n_22050;
assign n_22052 = ~x_142 &  n_22050;
assign n_22053 = ~n_22051 & ~n_22052;
assign n_22054 =  x_141 & ~n_21879;
assign n_22055 =  i_3 &  n_21879;
assign n_22056 = ~n_22054 & ~n_22055;
assign n_22057 =  x_141 & ~n_22056;
assign n_22058 = ~x_141 &  n_22056;
assign n_22059 = ~n_22057 & ~n_22058;
assign n_22060 =  x_140 & ~n_21879;
assign n_22061 =  i_2 &  n_21879;
assign n_22062 = ~n_22060 & ~n_22061;
assign n_22063 =  x_140 & ~n_22062;
assign n_22064 = ~x_140 &  n_22062;
assign n_22065 = ~n_22063 & ~n_22064;
assign n_22066 =  x_139 & ~n_21879;
assign n_22067 =  i_1 &  n_21879;
assign n_22068 = ~n_22066 & ~n_22067;
assign n_22069 =  x_139 & ~n_22068;
assign n_22070 = ~x_139 &  n_22068;
assign n_22071 = ~n_22069 & ~n_22070;
assign n_22072 =  n_1904 &  n_8254;
assign n_22073 =  x_138 & ~n_22072;
assign n_22074 =  i_32 &  n_22072;
assign n_22075 = ~n_22073 & ~n_22074;
assign n_22076 =  x_138 & ~n_22075;
assign n_22077 = ~x_138 &  n_22075;
assign n_22078 = ~n_22076 & ~n_22077;
assign n_22079 =  x_137 & ~n_22072;
assign n_22080 =  i_31 &  n_22072;
assign n_22081 = ~n_22079 & ~n_22080;
assign n_22082 =  x_137 & ~n_22081;
assign n_22083 = ~x_137 &  n_22081;
assign n_22084 = ~n_22082 & ~n_22083;
assign n_22085 =  x_136 & ~n_22072;
assign n_22086 =  i_30 &  n_22072;
assign n_22087 = ~n_22085 & ~n_22086;
assign n_22088 =  x_136 & ~n_22087;
assign n_22089 = ~x_136 &  n_22087;
assign n_22090 = ~n_22088 & ~n_22089;
assign n_22091 =  x_135 & ~n_22072;
assign n_22092 =  i_29 &  n_22072;
assign n_22093 = ~n_22091 & ~n_22092;
assign n_22094 =  x_135 & ~n_22093;
assign n_22095 = ~x_135 &  n_22093;
assign n_22096 = ~n_22094 & ~n_22095;
assign n_22097 =  x_134 & ~n_22072;
assign n_22098 =  i_28 &  n_22072;
assign n_22099 = ~n_22097 & ~n_22098;
assign n_22100 =  x_134 & ~n_22099;
assign n_22101 = ~x_134 &  n_22099;
assign n_22102 = ~n_22100 & ~n_22101;
assign n_22103 =  x_133 & ~n_22072;
assign n_22104 =  i_27 &  n_22072;
assign n_22105 = ~n_22103 & ~n_22104;
assign n_22106 =  x_133 & ~n_22105;
assign n_22107 = ~x_133 &  n_22105;
assign n_22108 = ~n_22106 & ~n_22107;
assign n_22109 =  x_132 & ~n_22072;
assign n_22110 =  i_26 &  n_22072;
assign n_22111 = ~n_22109 & ~n_22110;
assign n_22112 =  x_132 & ~n_22111;
assign n_22113 = ~x_132 &  n_22111;
assign n_22114 = ~n_22112 & ~n_22113;
assign n_22115 =  x_131 & ~n_22072;
assign n_22116 =  i_25 &  n_22072;
assign n_22117 = ~n_22115 & ~n_22116;
assign n_22118 =  x_131 & ~n_22117;
assign n_22119 = ~x_131 &  n_22117;
assign n_22120 = ~n_22118 & ~n_22119;
assign n_22121 =  x_130 & ~n_22072;
assign n_22122 =  i_24 &  n_22072;
assign n_22123 = ~n_22121 & ~n_22122;
assign n_22124 =  x_130 & ~n_22123;
assign n_22125 = ~x_130 &  n_22123;
assign n_22126 = ~n_22124 & ~n_22125;
assign n_22127 =  x_129 & ~n_22072;
assign n_22128 =  i_23 &  n_22072;
assign n_22129 = ~n_22127 & ~n_22128;
assign n_22130 =  x_129 & ~n_22129;
assign n_22131 = ~x_129 &  n_22129;
assign n_22132 = ~n_22130 & ~n_22131;
assign n_22133 =  x_128 & ~n_22072;
assign n_22134 =  i_22 &  n_22072;
assign n_22135 = ~n_22133 & ~n_22134;
assign n_22136 =  x_128 & ~n_22135;
assign n_22137 = ~x_128 &  n_22135;
assign n_22138 = ~n_22136 & ~n_22137;
assign n_22139 =  x_127 & ~n_22072;
assign n_22140 =  i_21 &  n_22072;
assign n_22141 = ~n_22139 & ~n_22140;
assign n_22142 =  x_127 & ~n_22141;
assign n_22143 = ~x_127 &  n_22141;
assign n_22144 = ~n_22142 & ~n_22143;
assign n_22145 =  x_126 & ~n_22072;
assign n_22146 =  i_20 &  n_22072;
assign n_22147 = ~n_22145 & ~n_22146;
assign n_22148 =  x_126 & ~n_22147;
assign n_22149 = ~x_126 &  n_22147;
assign n_22150 = ~n_22148 & ~n_22149;
assign n_22151 =  x_125 & ~n_22072;
assign n_22152 =  i_19 &  n_22072;
assign n_22153 = ~n_22151 & ~n_22152;
assign n_22154 =  x_125 & ~n_22153;
assign n_22155 = ~x_125 &  n_22153;
assign n_22156 = ~n_22154 & ~n_22155;
assign n_22157 =  x_124 & ~n_22072;
assign n_22158 =  i_18 &  n_22072;
assign n_22159 = ~n_22157 & ~n_22158;
assign n_22160 =  x_124 & ~n_22159;
assign n_22161 = ~x_124 &  n_22159;
assign n_22162 = ~n_22160 & ~n_22161;
assign n_22163 =  x_123 & ~n_22072;
assign n_22164 =  i_17 &  n_22072;
assign n_22165 = ~n_22163 & ~n_22164;
assign n_22166 =  x_123 & ~n_22165;
assign n_22167 = ~x_123 &  n_22165;
assign n_22168 = ~n_22166 & ~n_22167;
assign n_22169 =  x_122 & ~n_22072;
assign n_22170 =  i_16 &  n_22072;
assign n_22171 = ~n_22169 & ~n_22170;
assign n_22172 =  x_122 & ~n_22171;
assign n_22173 = ~x_122 &  n_22171;
assign n_22174 = ~n_22172 & ~n_22173;
assign n_22175 =  x_121 & ~n_22072;
assign n_22176 =  i_15 &  n_22072;
assign n_22177 = ~n_22175 & ~n_22176;
assign n_22178 =  x_121 & ~n_22177;
assign n_22179 = ~x_121 &  n_22177;
assign n_22180 = ~n_22178 & ~n_22179;
assign n_22181 =  x_120 & ~n_22072;
assign n_22182 =  i_14 &  n_22072;
assign n_22183 = ~n_22181 & ~n_22182;
assign n_22184 =  x_120 & ~n_22183;
assign n_22185 = ~x_120 &  n_22183;
assign n_22186 = ~n_22184 & ~n_22185;
assign n_22187 =  x_119 & ~n_22072;
assign n_22188 =  i_13 &  n_22072;
assign n_22189 = ~n_22187 & ~n_22188;
assign n_22190 =  x_119 & ~n_22189;
assign n_22191 = ~x_119 &  n_22189;
assign n_22192 = ~n_22190 & ~n_22191;
assign n_22193 =  x_118 & ~n_22072;
assign n_22194 =  i_12 &  n_22072;
assign n_22195 = ~n_22193 & ~n_22194;
assign n_22196 =  x_118 & ~n_22195;
assign n_22197 = ~x_118 &  n_22195;
assign n_22198 = ~n_22196 & ~n_22197;
assign n_22199 =  x_117 & ~n_22072;
assign n_22200 =  i_11 &  n_22072;
assign n_22201 = ~n_22199 & ~n_22200;
assign n_22202 =  x_117 & ~n_22201;
assign n_22203 = ~x_117 &  n_22201;
assign n_22204 = ~n_22202 & ~n_22203;
assign n_22205 =  x_116 & ~n_22072;
assign n_22206 =  i_10 &  n_22072;
assign n_22207 = ~n_22205 & ~n_22206;
assign n_22208 =  x_116 & ~n_22207;
assign n_22209 = ~x_116 &  n_22207;
assign n_22210 = ~n_22208 & ~n_22209;
assign n_22211 =  x_115 & ~n_22072;
assign n_22212 =  i_9 &  n_22072;
assign n_22213 = ~n_22211 & ~n_22212;
assign n_22214 =  x_115 & ~n_22213;
assign n_22215 = ~x_115 &  n_22213;
assign n_22216 = ~n_22214 & ~n_22215;
assign n_22217 =  x_114 & ~n_22072;
assign n_22218 =  i_8 &  n_22072;
assign n_22219 = ~n_22217 & ~n_22218;
assign n_22220 =  x_114 & ~n_22219;
assign n_22221 = ~x_114 &  n_22219;
assign n_22222 = ~n_22220 & ~n_22221;
assign n_22223 =  x_113 & ~n_22072;
assign n_22224 =  i_7 &  n_22072;
assign n_22225 = ~n_22223 & ~n_22224;
assign n_22226 =  x_113 & ~n_22225;
assign n_22227 = ~x_113 &  n_22225;
assign n_22228 = ~n_22226 & ~n_22227;
assign n_22229 =  x_112 & ~n_22072;
assign n_22230 =  i_6 &  n_22072;
assign n_22231 = ~n_22229 & ~n_22230;
assign n_22232 =  x_112 & ~n_22231;
assign n_22233 = ~x_112 &  n_22231;
assign n_22234 = ~n_22232 & ~n_22233;
assign n_22235 =  x_111 & ~n_22072;
assign n_22236 =  i_5 &  n_22072;
assign n_22237 = ~n_22235 & ~n_22236;
assign n_22238 =  x_111 & ~n_22237;
assign n_22239 = ~x_111 &  n_22237;
assign n_22240 = ~n_22238 & ~n_22239;
assign n_22241 =  x_110 & ~n_22072;
assign n_22242 =  i_4 &  n_22072;
assign n_22243 = ~n_22241 & ~n_22242;
assign n_22244 =  x_110 & ~n_22243;
assign n_22245 = ~x_110 &  n_22243;
assign n_22246 = ~n_22244 & ~n_22245;
assign n_22247 =  x_109 & ~n_22072;
assign n_22248 =  i_3 &  n_22072;
assign n_22249 = ~n_22247 & ~n_22248;
assign n_22250 =  x_109 & ~n_22249;
assign n_22251 = ~x_109 &  n_22249;
assign n_22252 = ~n_22250 & ~n_22251;
assign n_22253 =  x_108 & ~n_22072;
assign n_22254 =  i_2 &  n_22072;
assign n_22255 = ~n_22253 & ~n_22254;
assign n_22256 =  x_108 & ~n_22255;
assign n_22257 = ~x_108 &  n_22255;
assign n_22258 = ~n_22256 & ~n_22257;
assign n_22259 =  x_107 & ~n_22072;
assign n_22260 =  i_1 &  n_22072;
assign n_22261 = ~n_22259 & ~n_22260;
assign n_22262 =  x_107 & ~n_22261;
assign n_22263 = ~x_107 &  n_22261;
assign n_22264 = ~n_22262 & ~n_22263;
assign n_22265 =  n_586 &  n_2499;
assign n_22266 = ~x_39 &  n_22265;
assign n_22267 =  x_74 & ~n_22266;
assign n_22268 =  i_32 &  n_22266;
assign n_22269 = ~n_22267 & ~n_22268;
assign n_22270 =  x_74 & ~n_22269;
assign n_22271 = ~x_74 &  n_22269;
assign n_22272 = ~n_22270 & ~n_22271;
assign n_22273 =  x_73 & ~n_22266;
assign n_22274 =  i_31 &  n_22266;
assign n_22275 = ~n_22273 & ~n_22274;
assign n_22276 =  x_73 & ~n_22275;
assign n_22277 = ~x_73 &  n_22275;
assign n_22278 = ~n_22276 & ~n_22277;
assign n_22279 =  x_72 & ~n_22266;
assign n_22280 =  i_30 &  n_22266;
assign n_22281 = ~n_22279 & ~n_22280;
assign n_22282 =  x_72 & ~n_22281;
assign n_22283 = ~x_72 &  n_22281;
assign n_22284 = ~n_22282 & ~n_22283;
assign n_22285 =  x_71 & ~n_22266;
assign n_22286 =  i_29 &  n_22266;
assign n_22287 = ~n_22285 & ~n_22286;
assign n_22288 =  x_71 & ~n_22287;
assign n_22289 = ~x_71 &  n_22287;
assign n_22290 = ~n_22288 & ~n_22289;
assign n_22291 =  x_70 & ~n_22266;
assign n_22292 =  i_28 &  n_22266;
assign n_22293 = ~n_22291 & ~n_22292;
assign n_22294 =  x_70 & ~n_22293;
assign n_22295 = ~x_70 &  n_22293;
assign n_22296 = ~n_22294 & ~n_22295;
assign n_22297 =  x_69 & ~n_22266;
assign n_22298 =  i_27 &  n_22266;
assign n_22299 = ~n_22297 & ~n_22298;
assign n_22300 =  x_69 & ~n_22299;
assign n_22301 = ~x_69 &  n_22299;
assign n_22302 = ~n_22300 & ~n_22301;
assign n_22303 =  x_68 & ~n_22266;
assign n_22304 =  i_26 &  n_22266;
assign n_22305 = ~n_22303 & ~n_22304;
assign n_22306 =  x_68 & ~n_22305;
assign n_22307 = ~x_68 &  n_22305;
assign n_22308 = ~n_22306 & ~n_22307;
assign n_22309 =  x_67 & ~n_22266;
assign n_22310 =  i_25 &  n_22266;
assign n_22311 = ~n_22309 & ~n_22310;
assign n_22312 =  x_67 & ~n_22311;
assign n_22313 = ~x_67 &  n_22311;
assign n_22314 = ~n_22312 & ~n_22313;
assign n_22315 =  x_66 & ~n_22266;
assign n_22316 =  i_24 &  n_22266;
assign n_22317 = ~n_22315 & ~n_22316;
assign n_22318 =  x_66 & ~n_22317;
assign n_22319 = ~x_66 &  n_22317;
assign n_22320 = ~n_22318 & ~n_22319;
assign n_22321 =  x_65 & ~n_22266;
assign n_22322 =  i_23 &  n_22266;
assign n_22323 = ~n_22321 & ~n_22322;
assign n_22324 =  x_65 & ~n_22323;
assign n_22325 = ~x_65 &  n_22323;
assign n_22326 = ~n_22324 & ~n_22325;
assign n_22327 =  x_64 & ~n_22266;
assign n_22328 =  i_22 &  n_22266;
assign n_22329 = ~n_22327 & ~n_22328;
assign n_22330 =  x_64 & ~n_22329;
assign n_22331 = ~x_64 &  n_22329;
assign n_22332 = ~n_22330 & ~n_22331;
assign n_22333 =  x_63 & ~n_22266;
assign n_22334 =  i_21 &  n_22266;
assign n_22335 = ~n_22333 & ~n_22334;
assign n_22336 =  x_63 & ~n_22335;
assign n_22337 = ~x_63 &  n_22335;
assign n_22338 = ~n_22336 & ~n_22337;
assign n_22339 =  x_62 & ~n_22266;
assign n_22340 =  i_20 &  n_22266;
assign n_22341 = ~n_22339 & ~n_22340;
assign n_22342 =  x_62 & ~n_22341;
assign n_22343 = ~x_62 &  n_22341;
assign n_22344 = ~n_22342 & ~n_22343;
assign n_22345 =  n_586 &  n_18433;
assign n_22346 =  x_2858 & ~n_22345;
assign n_22347 =  i_32 &  n_22345;
assign n_22348 = ~n_22346 & ~n_22347;
assign n_22349 =  x_2858 & ~n_22348;
assign n_22350 = ~x_2858 &  n_22348;
assign n_22351 = ~n_22349 & ~n_22350;
assign n_22352 =  x_2857 & ~n_22345;
assign n_22353 =  i_31 &  n_22345;
assign n_22354 = ~n_22352 & ~n_22353;
assign n_22355 =  x_2857 & ~n_22354;
assign n_22356 = ~x_2857 &  n_22354;
assign n_22357 = ~n_22355 & ~n_22356;
assign n_22358 =  x_2856 & ~n_22345;
assign n_22359 =  i_30 &  n_22345;
assign n_22360 = ~n_22358 & ~n_22359;
assign n_22361 =  x_2856 & ~n_22360;
assign n_22362 = ~x_2856 &  n_22360;
assign n_22363 = ~n_22361 & ~n_22362;
assign n_22364 =  x_2855 & ~n_22345;
assign n_22365 =  i_29 &  n_22345;
assign n_22366 = ~n_22364 & ~n_22365;
assign n_22367 =  x_2855 & ~n_22366;
assign n_22368 = ~x_2855 &  n_22366;
assign n_22369 = ~n_22367 & ~n_22368;
assign n_22370 =  x_2854 & ~n_22345;
assign n_22371 =  i_28 &  n_22345;
assign n_22372 = ~n_22370 & ~n_22371;
assign n_22373 =  x_2854 & ~n_22372;
assign n_22374 = ~x_2854 &  n_22372;
assign n_22375 = ~n_22373 & ~n_22374;
assign n_22376 =  x_2853 & ~n_22345;
assign n_22377 =  i_27 &  n_22345;
assign n_22378 = ~n_22376 & ~n_22377;
assign n_22379 =  x_2853 & ~n_22378;
assign n_22380 = ~x_2853 &  n_22378;
assign n_22381 = ~n_22379 & ~n_22380;
assign n_22382 =  x_2852 & ~n_22345;
assign n_22383 =  i_26 &  n_22345;
assign n_22384 = ~n_22382 & ~n_22383;
assign n_22385 =  x_2852 & ~n_22384;
assign n_22386 = ~x_2852 &  n_22384;
assign n_22387 = ~n_22385 & ~n_22386;
assign n_22388 =  x_2851 & ~n_22345;
assign n_22389 =  i_25 &  n_22345;
assign n_22390 = ~n_22388 & ~n_22389;
assign n_22391 =  x_2851 & ~n_22390;
assign n_22392 = ~x_2851 &  n_22390;
assign n_22393 = ~n_22391 & ~n_22392;
assign n_22394 =  x_2850 & ~n_22345;
assign n_22395 =  i_24 &  n_22345;
assign n_22396 = ~n_22394 & ~n_22395;
assign n_22397 =  x_2850 & ~n_22396;
assign n_22398 = ~x_2850 &  n_22396;
assign n_22399 = ~n_22397 & ~n_22398;
assign n_22400 =  x_2849 & ~n_22345;
assign n_22401 =  i_23 &  n_22345;
assign n_22402 = ~n_22400 & ~n_22401;
assign n_22403 =  x_2849 & ~n_22402;
assign n_22404 = ~x_2849 &  n_22402;
assign n_22405 = ~n_22403 & ~n_22404;
assign n_22406 =  x_2848 & ~n_22345;
assign n_22407 =  i_22 &  n_22345;
assign n_22408 = ~n_22406 & ~n_22407;
assign n_22409 =  x_2848 & ~n_22408;
assign n_22410 = ~x_2848 &  n_22408;
assign n_22411 = ~n_22409 & ~n_22410;
assign n_22412 =  x_2847 & ~n_22345;
assign n_22413 =  i_21 &  n_22345;
assign n_22414 = ~n_22412 & ~n_22413;
assign n_22415 =  x_2847 & ~n_22414;
assign n_22416 = ~x_2847 &  n_22414;
assign n_22417 = ~n_22415 & ~n_22416;
assign n_22418 =  x_2846 & ~n_22345;
assign n_22419 =  i_20 &  n_22345;
assign n_22420 = ~n_22418 & ~n_22419;
assign n_22421 =  x_2846 & ~n_22420;
assign n_22422 = ~x_2846 &  n_22420;
assign n_22423 = ~n_22421 & ~n_22422;
assign n_22424 =  x_2845 & ~n_22345;
assign n_22425 =  i_19 &  n_22345;
assign n_22426 = ~n_22424 & ~n_22425;
assign n_22427 =  x_2845 & ~n_22426;
assign n_22428 = ~x_2845 &  n_22426;
assign n_22429 = ~n_22427 & ~n_22428;
assign n_22430 =  x_2844 & ~n_22345;
assign n_22431 =  i_18 &  n_22345;
assign n_22432 = ~n_22430 & ~n_22431;
assign n_22433 =  x_2844 & ~n_22432;
assign n_22434 = ~x_2844 &  n_22432;
assign n_22435 = ~n_22433 & ~n_22434;
assign n_22436 =  x_2843 & ~n_22345;
assign n_22437 =  i_17 &  n_22345;
assign n_22438 = ~n_22436 & ~n_22437;
assign n_22439 =  x_2843 & ~n_22438;
assign n_22440 = ~x_2843 &  n_22438;
assign n_22441 = ~n_22439 & ~n_22440;
assign n_22442 =  x_2842 & ~n_22345;
assign n_22443 =  i_16 &  n_22345;
assign n_22444 = ~n_22442 & ~n_22443;
assign n_22445 =  x_2842 & ~n_22444;
assign n_22446 = ~x_2842 &  n_22444;
assign n_22447 = ~n_22445 & ~n_22446;
assign n_22448 =  x_2841 & ~n_22345;
assign n_22449 =  i_15 &  n_22345;
assign n_22450 = ~n_22448 & ~n_22449;
assign n_22451 =  x_2841 & ~n_22450;
assign n_22452 = ~x_2841 &  n_22450;
assign n_22453 = ~n_22451 & ~n_22452;
assign n_22454 =  x_2840 & ~n_22345;
assign n_22455 =  i_14 &  n_22345;
assign n_22456 = ~n_22454 & ~n_22455;
assign n_22457 =  x_2840 & ~n_22456;
assign n_22458 = ~x_2840 &  n_22456;
assign n_22459 = ~n_22457 & ~n_22458;
assign n_22460 =  x_2839 & ~n_22345;
assign n_22461 =  i_13 &  n_22345;
assign n_22462 = ~n_22460 & ~n_22461;
assign n_22463 =  x_2839 & ~n_22462;
assign n_22464 = ~x_2839 &  n_22462;
assign n_22465 = ~n_22463 & ~n_22464;
assign n_22466 =  x_2838 & ~n_22345;
assign n_22467 =  i_12 &  n_22345;
assign n_22468 = ~n_22466 & ~n_22467;
assign n_22469 =  x_2838 & ~n_22468;
assign n_22470 = ~x_2838 &  n_22468;
assign n_22471 = ~n_22469 & ~n_22470;
assign n_22472 =  x_2837 & ~n_22345;
assign n_22473 =  i_11 &  n_22345;
assign n_22474 = ~n_22472 & ~n_22473;
assign n_22475 =  x_2837 & ~n_22474;
assign n_22476 = ~x_2837 &  n_22474;
assign n_22477 = ~n_22475 & ~n_22476;
assign n_22478 =  x_2836 & ~n_22345;
assign n_22479 =  i_10 &  n_22345;
assign n_22480 = ~n_22478 & ~n_22479;
assign n_22481 =  x_2836 & ~n_22480;
assign n_22482 = ~x_2836 &  n_22480;
assign n_22483 = ~n_22481 & ~n_22482;
assign n_22484 =  x_2835 & ~n_22345;
assign n_22485 =  i_9 &  n_22345;
assign n_22486 = ~n_22484 & ~n_22485;
assign n_22487 =  x_2835 & ~n_22486;
assign n_22488 = ~x_2835 &  n_22486;
assign n_22489 = ~n_22487 & ~n_22488;
assign n_22490 =  x_2834 & ~n_22345;
assign n_22491 =  i_8 &  n_22345;
assign n_22492 = ~n_22490 & ~n_22491;
assign n_22493 =  x_2834 & ~n_22492;
assign n_22494 = ~x_2834 &  n_22492;
assign n_22495 = ~n_22493 & ~n_22494;
assign n_22496 =  x_2833 & ~n_22345;
assign n_22497 =  i_7 &  n_22345;
assign n_22498 = ~n_22496 & ~n_22497;
assign n_22499 =  x_2833 & ~n_22498;
assign n_22500 = ~x_2833 &  n_22498;
assign n_22501 = ~n_22499 & ~n_22500;
assign n_22502 =  x_2832 & ~n_22345;
assign n_22503 =  i_6 &  n_22345;
assign n_22504 = ~n_22502 & ~n_22503;
assign n_22505 =  x_2832 & ~n_22504;
assign n_22506 = ~x_2832 &  n_22504;
assign n_22507 = ~n_22505 & ~n_22506;
assign n_22508 =  x_2831 & ~n_22345;
assign n_22509 =  i_5 &  n_22345;
assign n_22510 = ~n_22508 & ~n_22509;
assign n_22511 =  x_2831 & ~n_22510;
assign n_22512 = ~x_2831 &  n_22510;
assign n_22513 = ~n_22511 & ~n_22512;
assign n_22514 =  x_2830 & ~n_22345;
assign n_22515 =  i_4 &  n_22345;
assign n_22516 = ~n_22514 & ~n_22515;
assign n_22517 =  x_2830 & ~n_22516;
assign n_22518 = ~x_2830 &  n_22516;
assign n_22519 = ~n_22517 & ~n_22518;
assign n_22520 =  x_2829 & ~n_22345;
assign n_22521 =  i_3 &  n_22345;
assign n_22522 = ~n_22520 & ~n_22521;
assign n_22523 =  x_2829 & ~n_22522;
assign n_22524 = ~x_2829 &  n_22522;
assign n_22525 = ~n_22523 & ~n_22524;
assign n_22526 =  x_2828 & ~n_22345;
assign n_22527 =  i_2 &  n_22345;
assign n_22528 = ~n_22526 & ~n_22527;
assign n_22529 =  x_2828 & ~n_22528;
assign n_22530 = ~x_2828 &  n_22528;
assign n_22531 = ~n_22529 & ~n_22530;
assign n_22532 =  x_2827 & ~n_22345;
assign n_22533 =  i_1 &  n_22345;
assign n_22534 = ~n_22532 & ~n_22533;
assign n_22535 =  x_2827 & ~n_22534;
assign n_22536 = ~x_2827 &  n_22534;
assign n_22537 = ~n_22535 & ~n_22536;
assign n_22538 =  n_3664 &  n_1709;
assign n_22539 =  x_2826 & ~n_22538;
assign n_22540 =  i_32 &  n_22538;
assign n_22541 = ~n_22539 & ~n_22540;
assign n_22542 =  x_2826 & ~n_22541;
assign n_22543 = ~x_2826 &  n_22541;
assign n_22544 = ~n_22542 & ~n_22543;
assign n_22545 =  x_2825 & ~n_22538;
assign n_22546 =  i_31 &  n_22538;
assign n_22547 = ~n_22545 & ~n_22546;
assign n_22548 =  x_2825 & ~n_22547;
assign n_22549 = ~x_2825 &  n_22547;
assign n_22550 = ~n_22548 & ~n_22549;
assign n_22551 =  x_2824 & ~n_22538;
assign n_22552 =  i_30 &  n_22538;
assign n_22553 = ~n_22551 & ~n_22552;
assign n_22554 =  x_2824 & ~n_22553;
assign n_22555 = ~x_2824 &  n_22553;
assign n_22556 = ~n_22554 & ~n_22555;
assign n_22557 =  x_2823 & ~n_22538;
assign n_22558 =  i_29 &  n_22538;
assign n_22559 = ~n_22557 & ~n_22558;
assign n_22560 =  x_2823 & ~n_22559;
assign n_22561 = ~x_2823 &  n_22559;
assign n_22562 = ~n_22560 & ~n_22561;
assign n_22563 =  x_2822 & ~n_22538;
assign n_22564 =  i_28 &  n_22538;
assign n_22565 = ~n_22563 & ~n_22564;
assign n_22566 =  x_2822 & ~n_22565;
assign n_22567 = ~x_2822 &  n_22565;
assign n_22568 = ~n_22566 & ~n_22567;
assign n_22569 =  x_2821 & ~n_22538;
assign n_22570 =  i_27 &  n_22538;
assign n_22571 = ~n_22569 & ~n_22570;
assign n_22572 =  x_2821 & ~n_22571;
assign n_22573 = ~x_2821 &  n_22571;
assign n_22574 = ~n_22572 & ~n_22573;
assign n_22575 =  x_2820 & ~n_22538;
assign n_22576 =  i_26 &  n_22538;
assign n_22577 = ~n_22575 & ~n_22576;
assign n_22578 =  x_2820 & ~n_22577;
assign n_22579 = ~x_2820 &  n_22577;
assign n_22580 = ~n_22578 & ~n_22579;
assign n_22581 =  x_2819 & ~n_22538;
assign n_22582 =  i_25 &  n_22538;
assign n_22583 = ~n_22581 & ~n_22582;
assign n_22584 =  x_2819 & ~n_22583;
assign n_22585 = ~x_2819 &  n_22583;
assign n_22586 = ~n_22584 & ~n_22585;
assign n_22587 =  x_2818 & ~n_22538;
assign n_22588 =  i_24 &  n_22538;
assign n_22589 = ~n_22587 & ~n_22588;
assign n_22590 =  x_2818 & ~n_22589;
assign n_22591 = ~x_2818 &  n_22589;
assign n_22592 = ~n_22590 & ~n_22591;
assign n_22593 =  x_2817 & ~n_22538;
assign n_22594 =  i_23 &  n_22538;
assign n_22595 = ~n_22593 & ~n_22594;
assign n_22596 =  x_2817 & ~n_22595;
assign n_22597 = ~x_2817 &  n_22595;
assign n_22598 = ~n_22596 & ~n_22597;
assign n_22599 =  x_2816 & ~n_22538;
assign n_22600 =  i_22 &  n_22538;
assign n_22601 = ~n_22599 & ~n_22600;
assign n_22602 =  x_2816 & ~n_22601;
assign n_22603 = ~x_2816 &  n_22601;
assign n_22604 = ~n_22602 & ~n_22603;
assign n_22605 =  x_2815 & ~n_22538;
assign n_22606 =  i_21 &  n_22538;
assign n_22607 = ~n_22605 & ~n_22606;
assign n_22608 =  x_2815 & ~n_22607;
assign n_22609 = ~x_2815 &  n_22607;
assign n_22610 = ~n_22608 & ~n_22609;
assign n_22611 =  x_2814 & ~n_22538;
assign n_22612 =  i_20 &  n_22538;
assign n_22613 = ~n_22611 & ~n_22612;
assign n_22614 =  x_2814 & ~n_22613;
assign n_22615 = ~x_2814 &  n_22613;
assign n_22616 = ~n_22614 & ~n_22615;
assign n_22617 =  x_2813 & ~n_22538;
assign n_22618 =  i_19 &  n_22538;
assign n_22619 = ~n_22617 & ~n_22618;
assign n_22620 =  x_2813 & ~n_22619;
assign n_22621 = ~x_2813 &  n_22619;
assign n_22622 = ~n_22620 & ~n_22621;
assign n_22623 =  x_2812 & ~n_22538;
assign n_22624 =  i_18 &  n_22538;
assign n_22625 = ~n_22623 & ~n_22624;
assign n_22626 =  x_2812 & ~n_22625;
assign n_22627 = ~x_2812 &  n_22625;
assign n_22628 = ~n_22626 & ~n_22627;
assign n_22629 =  x_2811 & ~n_22538;
assign n_22630 =  i_17 &  n_22538;
assign n_22631 = ~n_22629 & ~n_22630;
assign n_22632 =  x_2811 & ~n_22631;
assign n_22633 = ~x_2811 &  n_22631;
assign n_22634 = ~n_22632 & ~n_22633;
assign n_22635 =  x_2810 & ~n_22538;
assign n_22636 =  i_16 &  n_22538;
assign n_22637 = ~n_22635 & ~n_22636;
assign n_22638 =  x_2810 & ~n_22637;
assign n_22639 = ~x_2810 &  n_22637;
assign n_22640 = ~n_22638 & ~n_22639;
assign n_22641 =  x_2809 & ~n_22538;
assign n_22642 =  i_15 &  n_22538;
assign n_22643 = ~n_22641 & ~n_22642;
assign n_22644 =  x_2809 & ~n_22643;
assign n_22645 = ~x_2809 &  n_22643;
assign n_22646 = ~n_22644 & ~n_22645;
assign n_22647 =  x_2808 & ~n_22538;
assign n_22648 =  i_14 &  n_22538;
assign n_22649 = ~n_22647 & ~n_22648;
assign n_22650 =  x_2808 & ~n_22649;
assign n_22651 = ~x_2808 &  n_22649;
assign n_22652 = ~n_22650 & ~n_22651;
assign n_22653 =  x_2807 & ~n_22538;
assign n_22654 =  i_13 &  n_22538;
assign n_22655 = ~n_22653 & ~n_22654;
assign n_22656 =  x_2807 & ~n_22655;
assign n_22657 = ~x_2807 &  n_22655;
assign n_22658 = ~n_22656 & ~n_22657;
assign n_22659 =  x_2806 & ~n_22538;
assign n_22660 =  i_12 &  n_22538;
assign n_22661 = ~n_22659 & ~n_22660;
assign n_22662 =  x_2806 & ~n_22661;
assign n_22663 = ~x_2806 &  n_22661;
assign n_22664 = ~n_22662 & ~n_22663;
assign n_22665 =  x_2805 & ~n_22538;
assign n_22666 =  i_11 &  n_22538;
assign n_22667 = ~n_22665 & ~n_22666;
assign n_22668 =  x_2805 & ~n_22667;
assign n_22669 = ~x_2805 &  n_22667;
assign n_22670 = ~n_22668 & ~n_22669;
assign n_22671 =  x_2804 & ~n_22538;
assign n_22672 =  i_10 &  n_22538;
assign n_22673 = ~n_22671 & ~n_22672;
assign n_22674 =  x_2804 & ~n_22673;
assign n_22675 = ~x_2804 &  n_22673;
assign n_22676 = ~n_22674 & ~n_22675;
assign n_22677 =  x_2803 & ~n_22538;
assign n_22678 =  i_9 &  n_22538;
assign n_22679 = ~n_22677 & ~n_22678;
assign n_22680 =  x_2803 & ~n_22679;
assign n_22681 = ~x_2803 &  n_22679;
assign n_22682 = ~n_22680 & ~n_22681;
assign n_22683 =  x_2802 & ~n_22538;
assign n_22684 =  i_8 &  n_22538;
assign n_22685 = ~n_22683 & ~n_22684;
assign n_22686 =  x_2802 & ~n_22685;
assign n_22687 = ~x_2802 &  n_22685;
assign n_22688 = ~n_22686 & ~n_22687;
assign n_22689 =  x_2801 & ~n_22538;
assign n_22690 =  i_7 &  n_22538;
assign n_22691 = ~n_22689 & ~n_22690;
assign n_22692 =  x_2801 & ~n_22691;
assign n_22693 = ~x_2801 &  n_22691;
assign n_22694 = ~n_22692 & ~n_22693;
assign n_22695 =  x_2800 & ~n_22538;
assign n_22696 =  i_6 &  n_22538;
assign n_22697 = ~n_22695 & ~n_22696;
assign n_22698 =  x_2800 & ~n_22697;
assign n_22699 = ~x_2800 &  n_22697;
assign n_22700 = ~n_22698 & ~n_22699;
assign n_22701 =  x_2799 & ~n_22538;
assign n_22702 =  i_5 &  n_22538;
assign n_22703 = ~n_22701 & ~n_22702;
assign n_22704 =  x_2799 & ~n_22703;
assign n_22705 = ~x_2799 &  n_22703;
assign n_22706 = ~n_22704 & ~n_22705;
assign n_22707 =  x_2798 & ~n_22538;
assign n_22708 =  i_4 &  n_22538;
assign n_22709 = ~n_22707 & ~n_22708;
assign n_22710 =  x_2798 & ~n_22709;
assign n_22711 = ~x_2798 &  n_22709;
assign n_22712 = ~n_22710 & ~n_22711;
assign n_22713 =  x_2797 & ~n_22538;
assign n_22714 =  i_3 &  n_22538;
assign n_22715 = ~n_22713 & ~n_22714;
assign n_22716 =  x_2797 & ~n_22715;
assign n_22717 = ~x_2797 &  n_22715;
assign n_22718 = ~n_22716 & ~n_22717;
assign n_22719 =  x_2796 & ~n_22538;
assign n_22720 =  i_2 &  n_22538;
assign n_22721 = ~n_22719 & ~n_22720;
assign n_22722 =  x_2796 & ~n_22721;
assign n_22723 = ~x_2796 &  n_22721;
assign n_22724 = ~n_22722 & ~n_22723;
assign n_22725 =  x_2795 & ~n_22538;
assign n_22726 =  i_1 &  n_22538;
assign n_22727 = ~n_22725 & ~n_22726;
assign n_22728 =  x_2795 & ~n_22727;
assign n_22729 = ~x_2795 &  n_22727;
assign n_22730 = ~n_22728 & ~n_22729;
assign n_22731 =  n_3858 &  n_1512;
assign n_22732 =  x_2794 & ~n_22731;
assign n_22733 =  i_32 &  n_22731;
assign n_22734 = ~n_22732 & ~n_22733;
assign n_22735 =  x_2794 & ~n_22734;
assign n_22736 = ~x_2794 &  n_22734;
assign n_22737 = ~n_22735 & ~n_22736;
assign n_22738 =  x_2793 & ~n_22731;
assign n_22739 =  i_31 &  n_22731;
assign n_22740 = ~n_22738 & ~n_22739;
assign n_22741 =  x_2793 & ~n_22740;
assign n_22742 = ~x_2793 &  n_22740;
assign n_22743 = ~n_22741 & ~n_22742;
assign n_22744 =  x_2792 & ~n_22731;
assign n_22745 =  i_30 &  n_22731;
assign n_22746 = ~n_22744 & ~n_22745;
assign n_22747 =  x_2792 & ~n_22746;
assign n_22748 = ~x_2792 &  n_22746;
assign n_22749 = ~n_22747 & ~n_22748;
assign n_22750 =  x_2791 & ~n_22731;
assign n_22751 =  i_29 &  n_22731;
assign n_22752 = ~n_22750 & ~n_22751;
assign n_22753 =  x_2791 & ~n_22752;
assign n_22754 = ~x_2791 &  n_22752;
assign n_22755 = ~n_22753 & ~n_22754;
assign n_22756 =  x_2790 & ~n_22731;
assign n_22757 =  i_28 &  n_22731;
assign n_22758 = ~n_22756 & ~n_22757;
assign n_22759 =  x_2790 & ~n_22758;
assign n_22760 = ~x_2790 &  n_22758;
assign n_22761 = ~n_22759 & ~n_22760;
assign n_22762 =  x_2789 & ~n_22731;
assign n_22763 =  i_27 &  n_22731;
assign n_22764 = ~n_22762 & ~n_22763;
assign n_22765 =  x_2789 & ~n_22764;
assign n_22766 = ~x_2789 &  n_22764;
assign n_22767 = ~n_22765 & ~n_22766;
assign n_22768 =  x_2788 & ~n_22731;
assign n_22769 =  i_26 &  n_22731;
assign n_22770 = ~n_22768 & ~n_22769;
assign n_22771 =  x_2788 & ~n_22770;
assign n_22772 = ~x_2788 &  n_22770;
assign n_22773 = ~n_22771 & ~n_22772;
assign n_22774 =  x_2787 & ~n_22731;
assign n_22775 =  i_25 &  n_22731;
assign n_22776 = ~n_22774 & ~n_22775;
assign n_22777 =  x_2787 & ~n_22776;
assign n_22778 = ~x_2787 &  n_22776;
assign n_22779 = ~n_22777 & ~n_22778;
assign n_22780 =  x_2786 & ~n_22731;
assign n_22781 =  i_24 &  n_22731;
assign n_22782 = ~n_22780 & ~n_22781;
assign n_22783 =  x_2786 & ~n_22782;
assign n_22784 = ~x_2786 &  n_22782;
assign n_22785 = ~n_22783 & ~n_22784;
assign n_22786 =  x_2785 & ~n_22731;
assign n_22787 =  i_23 &  n_22731;
assign n_22788 = ~n_22786 & ~n_22787;
assign n_22789 =  x_2785 & ~n_22788;
assign n_22790 = ~x_2785 &  n_22788;
assign n_22791 = ~n_22789 & ~n_22790;
assign n_22792 =  x_2784 & ~n_22731;
assign n_22793 =  i_22 &  n_22731;
assign n_22794 = ~n_22792 & ~n_22793;
assign n_22795 =  x_2784 & ~n_22794;
assign n_22796 = ~x_2784 &  n_22794;
assign n_22797 = ~n_22795 & ~n_22796;
assign n_22798 =  x_2783 & ~n_22731;
assign n_22799 =  i_21 &  n_22731;
assign n_22800 = ~n_22798 & ~n_22799;
assign n_22801 =  x_2783 & ~n_22800;
assign n_22802 = ~x_2783 &  n_22800;
assign n_22803 = ~n_22801 & ~n_22802;
assign n_22804 =  x_2782 & ~n_22731;
assign n_22805 =  i_20 &  n_22731;
assign n_22806 = ~n_22804 & ~n_22805;
assign n_22807 =  x_2782 & ~n_22806;
assign n_22808 = ~x_2782 &  n_22806;
assign n_22809 = ~n_22807 & ~n_22808;
assign n_22810 =  x_2781 & ~n_22731;
assign n_22811 =  i_19 &  n_22731;
assign n_22812 = ~n_22810 & ~n_22811;
assign n_22813 =  x_2781 & ~n_22812;
assign n_22814 = ~x_2781 &  n_22812;
assign n_22815 = ~n_22813 & ~n_22814;
assign n_22816 =  x_2780 & ~n_22731;
assign n_22817 =  i_18 &  n_22731;
assign n_22818 = ~n_22816 & ~n_22817;
assign n_22819 =  x_2780 & ~n_22818;
assign n_22820 = ~x_2780 &  n_22818;
assign n_22821 = ~n_22819 & ~n_22820;
assign n_22822 =  x_2779 & ~n_22731;
assign n_22823 =  i_17 &  n_22731;
assign n_22824 = ~n_22822 & ~n_22823;
assign n_22825 =  x_2779 & ~n_22824;
assign n_22826 = ~x_2779 &  n_22824;
assign n_22827 = ~n_22825 & ~n_22826;
assign n_22828 =  x_2778 & ~n_22731;
assign n_22829 =  i_16 &  n_22731;
assign n_22830 = ~n_22828 & ~n_22829;
assign n_22831 =  x_2778 & ~n_22830;
assign n_22832 = ~x_2778 &  n_22830;
assign n_22833 = ~n_22831 & ~n_22832;
assign n_22834 =  x_2777 & ~n_22731;
assign n_22835 =  i_15 &  n_22731;
assign n_22836 = ~n_22834 & ~n_22835;
assign n_22837 =  x_2777 & ~n_22836;
assign n_22838 = ~x_2777 &  n_22836;
assign n_22839 = ~n_22837 & ~n_22838;
assign n_22840 =  x_2776 & ~n_22731;
assign n_22841 =  i_14 &  n_22731;
assign n_22842 = ~n_22840 & ~n_22841;
assign n_22843 =  x_2776 & ~n_22842;
assign n_22844 = ~x_2776 &  n_22842;
assign n_22845 = ~n_22843 & ~n_22844;
assign n_22846 =  x_2775 & ~n_22731;
assign n_22847 =  i_13 &  n_22731;
assign n_22848 = ~n_22846 & ~n_22847;
assign n_22849 =  x_2775 & ~n_22848;
assign n_22850 = ~x_2775 &  n_22848;
assign n_22851 = ~n_22849 & ~n_22850;
assign n_22852 =  x_2774 & ~n_22731;
assign n_22853 =  i_12 &  n_22731;
assign n_22854 = ~n_22852 & ~n_22853;
assign n_22855 =  x_2774 & ~n_22854;
assign n_22856 = ~x_2774 &  n_22854;
assign n_22857 = ~n_22855 & ~n_22856;
assign n_22858 =  x_2773 & ~n_22731;
assign n_22859 =  i_11 &  n_22731;
assign n_22860 = ~n_22858 & ~n_22859;
assign n_22861 =  x_2773 & ~n_22860;
assign n_22862 = ~x_2773 &  n_22860;
assign n_22863 = ~n_22861 & ~n_22862;
assign n_22864 =  x_2772 & ~n_22731;
assign n_22865 =  i_10 &  n_22731;
assign n_22866 = ~n_22864 & ~n_22865;
assign n_22867 =  x_2772 & ~n_22866;
assign n_22868 = ~x_2772 &  n_22866;
assign n_22869 = ~n_22867 & ~n_22868;
assign n_22870 =  x_2771 & ~n_22731;
assign n_22871 =  i_9 &  n_22731;
assign n_22872 = ~n_22870 & ~n_22871;
assign n_22873 =  x_2771 & ~n_22872;
assign n_22874 = ~x_2771 &  n_22872;
assign n_22875 = ~n_22873 & ~n_22874;
assign n_22876 =  x_2770 & ~n_22731;
assign n_22877 =  i_8 &  n_22731;
assign n_22878 = ~n_22876 & ~n_22877;
assign n_22879 =  x_2770 & ~n_22878;
assign n_22880 = ~x_2770 &  n_22878;
assign n_22881 = ~n_22879 & ~n_22880;
assign n_22882 =  x_2769 & ~n_22731;
assign n_22883 =  i_7 &  n_22731;
assign n_22884 = ~n_22882 & ~n_22883;
assign n_22885 =  x_2769 & ~n_22884;
assign n_22886 = ~x_2769 &  n_22884;
assign n_22887 = ~n_22885 & ~n_22886;
assign n_22888 =  x_2768 & ~n_22731;
assign n_22889 =  i_6 &  n_22731;
assign n_22890 = ~n_22888 & ~n_22889;
assign n_22891 =  x_2768 & ~n_22890;
assign n_22892 = ~x_2768 &  n_22890;
assign n_22893 = ~n_22891 & ~n_22892;
assign n_22894 =  x_2767 & ~n_22731;
assign n_22895 =  i_5 &  n_22731;
assign n_22896 = ~n_22894 & ~n_22895;
assign n_22897 =  x_2767 & ~n_22896;
assign n_22898 = ~x_2767 &  n_22896;
assign n_22899 = ~n_22897 & ~n_22898;
assign n_22900 =  x_2766 & ~n_22731;
assign n_22901 =  i_4 &  n_22731;
assign n_22902 = ~n_22900 & ~n_22901;
assign n_22903 =  x_2766 & ~n_22902;
assign n_22904 = ~x_2766 &  n_22902;
assign n_22905 = ~n_22903 & ~n_22904;
assign n_22906 =  x_2765 & ~n_22731;
assign n_22907 =  i_3 &  n_22731;
assign n_22908 = ~n_22906 & ~n_22907;
assign n_22909 =  x_2765 & ~n_22908;
assign n_22910 = ~x_2765 &  n_22908;
assign n_22911 = ~n_22909 & ~n_22910;
assign n_22912 =  x_2764 & ~n_22731;
assign n_22913 =  i_2 &  n_22731;
assign n_22914 = ~n_22912 & ~n_22913;
assign n_22915 =  x_2764 & ~n_22914;
assign n_22916 = ~x_2764 &  n_22914;
assign n_22917 = ~n_22915 & ~n_22916;
assign n_22918 =  x_2763 & ~n_22731;
assign n_22919 =  i_1 &  n_22731;
assign n_22920 = ~n_22918 & ~n_22919;
assign n_22921 =  x_2763 & ~n_22920;
assign n_22922 = ~x_2763 &  n_22920;
assign n_22923 = ~n_22921 & ~n_22922;
assign n_22924 =  n_3664 &  n_6532;
assign n_22925 =  x_2762 & ~n_22924;
assign n_22926 =  i_32 &  n_22924;
assign n_22927 = ~n_22925 & ~n_22926;
assign n_22928 =  x_2762 & ~n_22927;
assign n_22929 = ~x_2762 &  n_22927;
assign n_22930 = ~n_22928 & ~n_22929;
assign n_22931 =  x_2761 & ~n_22924;
assign n_22932 =  i_31 &  n_22924;
assign n_22933 = ~n_22931 & ~n_22932;
assign n_22934 =  x_2761 & ~n_22933;
assign n_22935 = ~x_2761 &  n_22933;
assign n_22936 = ~n_22934 & ~n_22935;
assign n_22937 =  x_2760 & ~n_22924;
assign n_22938 =  i_30 &  n_22924;
assign n_22939 = ~n_22937 & ~n_22938;
assign n_22940 =  x_2760 & ~n_22939;
assign n_22941 = ~x_2760 &  n_22939;
assign n_22942 = ~n_22940 & ~n_22941;
assign n_22943 =  x_2759 & ~n_22924;
assign n_22944 =  i_29 &  n_22924;
assign n_22945 = ~n_22943 & ~n_22944;
assign n_22946 =  x_2759 & ~n_22945;
assign n_22947 = ~x_2759 &  n_22945;
assign n_22948 = ~n_22946 & ~n_22947;
assign n_22949 =  x_2758 & ~n_22924;
assign n_22950 =  i_28 &  n_22924;
assign n_22951 = ~n_22949 & ~n_22950;
assign n_22952 =  x_2758 & ~n_22951;
assign n_22953 = ~x_2758 &  n_22951;
assign n_22954 = ~n_22952 & ~n_22953;
assign n_22955 =  x_2757 & ~n_22924;
assign n_22956 =  i_27 &  n_22924;
assign n_22957 = ~n_22955 & ~n_22956;
assign n_22958 =  x_2757 & ~n_22957;
assign n_22959 = ~x_2757 &  n_22957;
assign n_22960 = ~n_22958 & ~n_22959;
assign n_22961 =  x_2756 & ~n_22924;
assign n_22962 =  i_26 &  n_22924;
assign n_22963 = ~n_22961 & ~n_22962;
assign n_22964 =  x_2756 & ~n_22963;
assign n_22965 = ~x_2756 &  n_22963;
assign n_22966 = ~n_22964 & ~n_22965;
assign n_22967 =  x_2755 & ~n_22924;
assign n_22968 =  i_25 &  n_22924;
assign n_22969 = ~n_22967 & ~n_22968;
assign n_22970 =  x_2755 & ~n_22969;
assign n_22971 = ~x_2755 &  n_22969;
assign n_22972 = ~n_22970 & ~n_22971;
assign n_22973 =  x_2754 & ~n_22924;
assign n_22974 =  i_24 &  n_22924;
assign n_22975 = ~n_22973 & ~n_22974;
assign n_22976 =  x_2754 & ~n_22975;
assign n_22977 = ~x_2754 &  n_22975;
assign n_22978 = ~n_22976 & ~n_22977;
assign n_22979 =  x_2753 & ~n_22924;
assign n_22980 =  i_23 &  n_22924;
assign n_22981 = ~n_22979 & ~n_22980;
assign n_22982 =  x_2753 & ~n_22981;
assign n_22983 = ~x_2753 &  n_22981;
assign n_22984 = ~n_22982 & ~n_22983;
assign n_22985 =  x_2752 & ~n_22924;
assign n_22986 =  i_22 &  n_22924;
assign n_22987 = ~n_22985 & ~n_22986;
assign n_22988 =  x_2752 & ~n_22987;
assign n_22989 = ~x_2752 &  n_22987;
assign n_22990 = ~n_22988 & ~n_22989;
assign n_22991 =  x_2751 & ~n_22924;
assign n_22992 =  i_21 &  n_22924;
assign n_22993 = ~n_22991 & ~n_22992;
assign n_22994 =  x_2751 & ~n_22993;
assign n_22995 = ~x_2751 &  n_22993;
assign n_22996 = ~n_22994 & ~n_22995;
assign n_22997 =  x_2750 & ~n_22924;
assign n_22998 =  i_20 &  n_22924;
assign n_22999 = ~n_22997 & ~n_22998;
assign n_23000 =  x_2750 & ~n_22999;
assign n_23001 = ~x_2750 &  n_22999;
assign n_23002 = ~n_23000 & ~n_23001;
assign n_23003 =  x_2749 & ~n_22924;
assign n_23004 =  i_19 &  n_22924;
assign n_23005 = ~n_23003 & ~n_23004;
assign n_23006 =  x_2749 & ~n_23005;
assign n_23007 = ~x_2749 &  n_23005;
assign n_23008 = ~n_23006 & ~n_23007;
assign n_23009 =  x_2748 & ~n_22924;
assign n_23010 =  i_18 &  n_22924;
assign n_23011 = ~n_23009 & ~n_23010;
assign n_23012 =  x_2748 & ~n_23011;
assign n_23013 = ~x_2748 &  n_23011;
assign n_23014 = ~n_23012 & ~n_23013;
assign n_23015 =  x_2747 & ~n_22924;
assign n_23016 =  i_17 &  n_22924;
assign n_23017 = ~n_23015 & ~n_23016;
assign n_23018 =  x_2747 & ~n_23017;
assign n_23019 = ~x_2747 &  n_23017;
assign n_23020 = ~n_23018 & ~n_23019;
assign n_23021 =  x_2746 & ~n_22924;
assign n_23022 =  i_16 &  n_22924;
assign n_23023 = ~n_23021 & ~n_23022;
assign n_23024 =  x_2746 & ~n_23023;
assign n_23025 = ~x_2746 &  n_23023;
assign n_23026 = ~n_23024 & ~n_23025;
assign n_23027 =  x_2745 & ~n_22924;
assign n_23028 =  i_15 &  n_22924;
assign n_23029 = ~n_23027 & ~n_23028;
assign n_23030 =  x_2745 & ~n_23029;
assign n_23031 = ~x_2745 &  n_23029;
assign n_23032 = ~n_23030 & ~n_23031;
assign n_23033 =  x_2744 & ~n_22924;
assign n_23034 =  i_14 &  n_22924;
assign n_23035 = ~n_23033 & ~n_23034;
assign n_23036 =  x_2744 & ~n_23035;
assign n_23037 = ~x_2744 &  n_23035;
assign n_23038 = ~n_23036 & ~n_23037;
assign n_23039 =  x_2743 & ~n_22924;
assign n_23040 =  i_13 &  n_22924;
assign n_23041 = ~n_23039 & ~n_23040;
assign n_23042 =  x_2743 & ~n_23041;
assign n_23043 = ~x_2743 &  n_23041;
assign n_23044 = ~n_23042 & ~n_23043;
assign n_23045 =  x_2742 & ~n_22924;
assign n_23046 =  i_12 &  n_22924;
assign n_23047 = ~n_23045 & ~n_23046;
assign n_23048 =  x_2742 & ~n_23047;
assign n_23049 = ~x_2742 &  n_23047;
assign n_23050 = ~n_23048 & ~n_23049;
assign n_23051 =  x_2741 & ~n_22924;
assign n_23052 =  i_11 &  n_22924;
assign n_23053 = ~n_23051 & ~n_23052;
assign n_23054 =  x_2741 & ~n_23053;
assign n_23055 = ~x_2741 &  n_23053;
assign n_23056 = ~n_23054 & ~n_23055;
assign n_23057 =  x_2740 & ~n_22924;
assign n_23058 =  i_10 &  n_22924;
assign n_23059 = ~n_23057 & ~n_23058;
assign n_23060 =  x_2740 & ~n_23059;
assign n_23061 = ~x_2740 &  n_23059;
assign n_23062 = ~n_23060 & ~n_23061;
assign n_23063 =  x_2739 & ~n_22924;
assign n_23064 =  i_9 &  n_22924;
assign n_23065 = ~n_23063 & ~n_23064;
assign n_23066 =  x_2739 & ~n_23065;
assign n_23067 = ~x_2739 &  n_23065;
assign n_23068 = ~n_23066 & ~n_23067;
assign n_23069 =  x_2738 & ~n_22924;
assign n_23070 =  i_8 &  n_22924;
assign n_23071 = ~n_23069 & ~n_23070;
assign n_23072 =  x_2738 & ~n_23071;
assign n_23073 = ~x_2738 &  n_23071;
assign n_23074 = ~n_23072 & ~n_23073;
assign n_23075 =  x_2737 & ~n_22924;
assign n_23076 =  i_7 &  n_22924;
assign n_23077 = ~n_23075 & ~n_23076;
assign n_23078 =  x_2737 & ~n_23077;
assign n_23079 = ~x_2737 &  n_23077;
assign n_23080 = ~n_23078 & ~n_23079;
assign n_23081 =  x_2736 & ~n_22924;
assign n_23082 =  i_6 &  n_22924;
assign n_23083 = ~n_23081 & ~n_23082;
assign n_23084 =  x_2736 & ~n_23083;
assign n_23085 = ~x_2736 &  n_23083;
assign n_23086 = ~n_23084 & ~n_23085;
assign n_23087 =  x_2735 & ~n_22924;
assign n_23088 =  i_5 &  n_22924;
assign n_23089 = ~n_23087 & ~n_23088;
assign n_23090 =  x_2735 & ~n_23089;
assign n_23091 = ~x_2735 &  n_23089;
assign n_23092 = ~n_23090 & ~n_23091;
assign n_23093 =  x_2734 & ~n_22924;
assign n_23094 =  i_4 &  n_22924;
assign n_23095 = ~n_23093 & ~n_23094;
assign n_23096 =  x_2734 & ~n_23095;
assign n_23097 = ~x_2734 &  n_23095;
assign n_23098 = ~n_23096 & ~n_23097;
assign n_23099 =  x_2733 & ~n_22924;
assign n_23100 =  i_3 &  n_22924;
assign n_23101 = ~n_23099 & ~n_23100;
assign n_23102 =  x_2733 & ~n_23101;
assign n_23103 = ~x_2733 &  n_23101;
assign n_23104 = ~n_23102 & ~n_23103;
assign n_23105 =  x_2732 & ~n_22924;
assign n_23106 =  i_2 &  n_22924;
assign n_23107 = ~n_23105 & ~n_23106;
assign n_23108 =  x_2732 & ~n_23107;
assign n_23109 = ~x_2732 &  n_23107;
assign n_23110 = ~n_23108 & ~n_23109;
assign n_23111 =  x_2731 & ~n_22924;
assign n_23112 =  i_1 &  n_22924;
assign n_23113 = ~n_23111 & ~n_23112;
assign n_23114 =  x_2731 & ~n_23113;
assign n_23115 = ~x_2731 &  n_23113;
assign n_23116 = ~n_23114 & ~n_23115;
assign n_23117 =  n_3 &  n_390;
assign n_23118 =  x_2730 & ~n_23117;
assign n_23119 =  i_32 &  n_23117;
assign n_23120 = ~n_23118 & ~n_23119;
assign n_23121 =  x_2730 & ~n_23120;
assign n_23122 = ~x_2730 &  n_23120;
assign n_23123 = ~n_23121 & ~n_23122;
assign n_23124 =  x_2729 & ~n_23117;
assign n_23125 =  i_31 &  n_23117;
assign n_23126 = ~n_23124 & ~n_23125;
assign n_23127 =  x_2729 & ~n_23126;
assign n_23128 = ~x_2729 &  n_23126;
assign n_23129 = ~n_23127 & ~n_23128;
assign n_23130 =  x_2728 & ~n_23117;
assign n_23131 =  i_30 &  n_23117;
assign n_23132 = ~n_23130 & ~n_23131;
assign n_23133 =  x_2728 & ~n_23132;
assign n_23134 = ~x_2728 &  n_23132;
assign n_23135 = ~n_23133 & ~n_23134;
assign n_23136 =  x_2727 & ~n_23117;
assign n_23137 =  i_29 &  n_23117;
assign n_23138 = ~n_23136 & ~n_23137;
assign n_23139 =  x_2727 & ~n_23138;
assign n_23140 = ~x_2727 &  n_23138;
assign n_23141 = ~n_23139 & ~n_23140;
assign n_23142 =  x_2726 & ~n_23117;
assign n_23143 =  i_28 &  n_23117;
assign n_23144 = ~n_23142 & ~n_23143;
assign n_23145 =  x_2726 & ~n_23144;
assign n_23146 = ~x_2726 &  n_23144;
assign n_23147 = ~n_23145 & ~n_23146;
assign n_23148 =  x_2725 & ~n_23117;
assign n_23149 =  i_27 &  n_23117;
assign n_23150 = ~n_23148 & ~n_23149;
assign n_23151 =  x_2725 & ~n_23150;
assign n_23152 = ~x_2725 &  n_23150;
assign n_23153 = ~n_23151 & ~n_23152;
assign n_23154 =  x_2724 & ~n_23117;
assign n_23155 =  i_26 &  n_23117;
assign n_23156 = ~n_23154 & ~n_23155;
assign n_23157 =  x_2724 & ~n_23156;
assign n_23158 = ~x_2724 &  n_23156;
assign n_23159 = ~n_23157 & ~n_23158;
assign n_23160 =  x_2723 & ~n_23117;
assign n_23161 =  i_25 &  n_23117;
assign n_23162 = ~n_23160 & ~n_23161;
assign n_23163 =  x_2723 & ~n_23162;
assign n_23164 = ~x_2723 &  n_23162;
assign n_23165 = ~n_23163 & ~n_23164;
assign n_23166 =  x_2722 & ~n_23117;
assign n_23167 =  i_24 &  n_23117;
assign n_23168 = ~n_23166 & ~n_23167;
assign n_23169 =  x_2722 & ~n_23168;
assign n_23170 = ~x_2722 &  n_23168;
assign n_23171 = ~n_23169 & ~n_23170;
assign n_23172 =  x_2721 & ~n_23117;
assign n_23173 =  i_23 &  n_23117;
assign n_23174 = ~n_23172 & ~n_23173;
assign n_23175 =  x_2721 & ~n_23174;
assign n_23176 = ~x_2721 &  n_23174;
assign n_23177 = ~n_23175 & ~n_23176;
assign n_23178 =  x_2720 & ~n_23117;
assign n_23179 =  i_22 &  n_23117;
assign n_23180 = ~n_23178 & ~n_23179;
assign n_23181 =  x_2720 & ~n_23180;
assign n_23182 = ~x_2720 &  n_23180;
assign n_23183 = ~n_23181 & ~n_23182;
assign n_23184 =  x_2719 & ~n_23117;
assign n_23185 =  i_21 &  n_23117;
assign n_23186 = ~n_23184 & ~n_23185;
assign n_23187 =  x_2719 & ~n_23186;
assign n_23188 = ~x_2719 &  n_23186;
assign n_23189 = ~n_23187 & ~n_23188;
assign n_23190 =  x_2718 & ~n_23117;
assign n_23191 =  i_20 &  n_23117;
assign n_23192 = ~n_23190 & ~n_23191;
assign n_23193 =  x_2718 & ~n_23192;
assign n_23194 = ~x_2718 &  n_23192;
assign n_23195 = ~n_23193 & ~n_23194;
assign n_23196 =  x_2717 & ~n_23117;
assign n_23197 =  i_19 &  n_23117;
assign n_23198 = ~n_23196 & ~n_23197;
assign n_23199 =  x_2717 & ~n_23198;
assign n_23200 = ~x_2717 &  n_23198;
assign n_23201 = ~n_23199 & ~n_23200;
assign n_23202 =  x_2716 & ~n_23117;
assign n_23203 =  i_18 &  n_23117;
assign n_23204 = ~n_23202 & ~n_23203;
assign n_23205 =  x_2716 & ~n_23204;
assign n_23206 = ~x_2716 &  n_23204;
assign n_23207 = ~n_23205 & ~n_23206;
assign n_23208 =  x_2715 & ~n_23117;
assign n_23209 =  i_17 &  n_23117;
assign n_23210 = ~n_23208 & ~n_23209;
assign n_23211 =  x_2715 & ~n_23210;
assign n_23212 = ~x_2715 &  n_23210;
assign n_23213 = ~n_23211 & ~n_23212;
assign n_23214 =  x_2714 & ~n_23117;
assign n_23215 =  i_16 &  n_23117;
assign n_23216 = ~n_23214 & ~n_23215;
assign n_23217 =  x_2714 & ~n_23216;
assign n_23218 = ~x_2714 &  n_23216;
assign n_23219 = ~n_23217 & ~n_23218;
assign n_23220 =  x_2713 & ~n_23117;
assign n_23221 =  i_15 &  n_23117;
assign n_23222 = ~n_23220 & ~n_23221;
assign n_23223 =  x_2713 & ~n_23222;
assign n_23224 = ~x_2713 &  n_23222;
assign n_23225 = ~n_23223 & ~n_23224;
assign n_23226 =  x_2712 & ~n_23117;
assign n_23227 =  i_14 &  n_23117;
assign n_23228 = ~n_23226 & ~n_23227;
assign n_23229 =  x_2712 & ~n_23228;
assign n_23230 = ~x_2712 &  n_23228;
assign n_23231 = ~n_23229 & ~n_23230;
assign n_23232 =  x_2711 & ~n_23117;
assign n_23233 =  i_13 &  n_23117;
assign n_23234 = ~n_23232 & ~n_23233;
assign n_23235 =  x_2711 & ~n_23234;
assign n_23236 = ~x_2711 &  n_23234;
assign n_23237 = ~n_23235 & ~n_23236;
assign n_23238 =  x_2710 & ~n_23117;
assign n_23239 =  i_12 &  n_23117;
assign n_23240 = ~n_23238 & ~n_23239;
assign n_23241 =  x_2710 & ~n_23240;
assign n_23242 = ~x_2710 &  n_23240;
assign n_23243 = ~n_23241 & ~n_23242;
assign n_23244 =  x_2709 & ~n_23117;
assign n_23245 =  i_11 &  n_23117;
assign n_23246 = ~n_23244 & ~n_23245;
assign n_23247 =  x_2709 & ~n_23246;
assign n_23248 = ~x_2709 &  n_23246;
assign n_23249 = ~n_23247 & ~n_23248;
assign n_23250 =  x_2708 & ~n_23117;
assign n_23251 =  i_10 &  n_23117;
assign n_23252 = ~n_23250 & ~n_23251;
assign n_23253 =  x_2708 & ~n_23252;
assign n_23254 = ~x_2708 &  n_23252;
assign n_23255 = ~n_23253 & ~n_23254;
assign n_23256 =  x_2707 & ~n_23117;
assign n_23257 =  i_9 &  n_23117;
assign n_23258 = ~n_23256 & ~n_23257;
assign n_23259 =  x_2707 & ~n_23258;
assign n_23260 = ~x_2707 &  n_23258;
assign n_23261 = ~n_23259 & ~n_23260;
assign n_23262 =  x_2706 & ~n_23117;
assign n_23263 =  i_8 &  n_23117;
assign n_23264 = ~n_23262 & ~n_23263;
assign n_23265 =  x_2706 & ~n_23264;
assign n_23266 = ~x_2706 &  n_23264;
assign n_23267 = ~n_23265 & ~n_23266;
assign n_23268 =  x_2705 & ~n_23117;
assign n_23269 =  i_7 &  n_23117;
assign n_23270 = ~n_23268 & ~n_23269;
assign n_23271 =  x_2705 & ~n_23270;
assign n_23272 = ~x_2705 &  n_23270;
assign n_23273 = ~n_23271 & ~n_23272;
assign n_23274 =  x_2704 & ~n_23117;
assign n_23275 =  i_6 &  n_23117;
assign n_23276 = ~n_23274 & ~n_23275;
assign n_23277 =  x_2704 & ~n_23276;
assign n_23278 = ~x_2704 &  n_23276;
assign n_23279 = ~n_23277 & ~n_23278;
assign n_23280 =  x_2703 & ~n_23117;
assign n_23281 =  i_5 &  n_23117;
assign n_23282 = ~n_23280 & ~n_23281;
assign n_23283 =  x_2703 & ~n_23282;
assign n_23284 = ~x_2703 &  n_23282;
assign n_23285 = ~n_23283 & ~n_23284;
assign n_23286 =  x_2702 & ~n_23117;
assign n_23287 =  i_4 &  n_23117;
assign n_23288 = ~n_23286 & ~n_23287;
assign n_23289 =  x_2702 & ~n_23288;
assign n_23290 = ~x_2702 &  n_23288;
assign n_23291 = ~n_23289 & ~n_23290;
assign n_23292 =  x_2701 & ~n_23117;
assign n_23293 =  i_3 &  n_23117;
assign n_23294 = ~n_23292 & ~n_23293;
assign n_23295 =  x_2701 & ~n_23294;
assign n_23296 = ~x_2701 &  n_23294;
assign n_23297 = ~n_23295 & ~n_23296;
assign n_23298 =  x_2700 & ~n_23117;
assign n_23299 =  i_2 &  n_23117;
assign n_23300 = ~n_23298 & ~n_23299;
assign n_23301 =  x_2700 & ~n_23300;
assign n_23302 = ~x_2700 &  n_23300;
assign n_23303 = ~n_23301 & ~n_23302;
assign n_23304 =  x_2699 & ~n_23117;
assign n_23305 =  i_1 &  n_23117;
assign n_23306 = ~n_23304 & ~n_23305;
assign n_23307 =  x_2699 & ~n_23306;
assign n_23308 = ~x_2699 &  n_23306;
assign n_23309 = ~n_23307 & ~n_23308;
assign n_23310 =  n_1315 &  n_10518;
assign n_23311 =  x_2698 & ~n_23310;
assign n_23312 =  i_32 &  n_23310;
assign n_23313 = ~n_23311 & ~n_23312;
assign n_23314 =  x_2698 & ~n_23313;
assign n_23315 = ~x_2698 &  n_23313;
assign n_23316 = ~n_23314 & ~n_23315;
assign n_23317 =  x_2697 & ~n_23310;
assign n_23318 =  i_31 &  n_23310;
assign n_23319 = ~n_23317 & ~n_23318;
assign n_23320 =  x_2697 & ~n_23319;
assign n_23321 = ~x_2697 &  n_23319;
assign n_23322 = ~n_23320 & ~n_23321;
assign n_23323 =  x_2696 & ~n_23310;
assign n_23324 =  i_30 &  n_23310;
assign n_23325 = ~n_23323 & ~n_23324;
assign n_23326 =  x_2696 & ~n_23325;
assign n_23327 = ~x_2696 &  n_23325;
assign n_23328 = ~n_23326 & ~n_23327;
assign n_23329 =  x_2695 & ~n_23310;
assign n_23330 =  i_29 &  n_23310;
assign n_23331 = ~n_23329 & ~n_23330;
assign n_23332 =  x_2695 & ~n_23331;
assign n_23333 = ~x_2695 &  n_23331;
assign n_23334 = ~n_23332 & ~n_23333;
assign n_23335 =  x_2694 & ~n_23310;
assign n_23336 =  i_28 &  n_23310;
assign n_23337 = ~n_23335 & ~n_23336;
assign n_23338 =  x_2694 & ~n_23337;
assign n_23339 = ~x_2694 &  n_23337;
assign n_23340 = ~n_23338 & ~n_23339;
assign n_23341 =  x_2693 & ~n_23310;
assign n_23342 =  i_27 &  n_23310;
assign n_23343 = ~n_23341 & ~n_23342;
assign n_23344 =  x_2693 & ~n_23343;
assign n_23345 = ~x_2693 &  n_23343;
assign n_23346 = ~n_23344 & ~n_23345;
assign n_23347 =  x_2692 & ~n_23310;
assign n_23348 =  i_26 &  n_23310;
assign n_23349 = ~n_23347 & ~n_23348;
assign n_23350 =  x_2692 & ~n_23349;
assign n_23351 = ~x_2692 &  n_23349;
assign n_23352 = ~n_23350 & ~n_23351;
assign n_23353 =  x_2691 & ~n_23310;
assign n_23354 =  i_25 &  n_23310;
assign n_23355 = ~n_23353 & ~n_23354;
assign n_23356 =  x_2691 & ~n_23355;
assign n_23357 = ~x_2691 &  n_23355;
assign n_23358 = ~n_23356 & ~n_23357;
assign n_23359 =  x_2690 & ~n_23310;
assign n_23360 =  i_24 &  n_23310;
assign n_23361 = ~n_23359 & ~n_23360;
assign n_23362 =  x_2690 & ~n_23361;
assign n_23363 = ~x_2690 &  n_23361;
assign n_23364 = ~n_23362 & ~n_23363;
assign n_23365 =  x_2689 & ~n_23310;
assign n_23366 =  i_23 &  n_23310;
assign n_23367 = ~n_23365 & ~n_23366;
assign n_23368 =  x_2689 & ~n_23367;
assign n_23369 = ~x_2689 &  n_23367;
assign n_23370 = ~n_23368 & ~n_23369;
assign n_23371 =  x_2688 & ~n_23310;
assign n_23372 =  i_22 &  n_23310;
assign n_23373 = ~n_23371 & ~n_23372;
assign n_23374 =  x_2688 & ~n_23373;
assign n_23375 = ~x_2688 &  n_23373;
assign n_23376 = ~n_23374 & ~n_23375;
assign n_23377 =  x_2687 & ~n_23310;
assign n_23378 =  i_21 &  n_23310;
assign n_23379 = ~n_23377 & ~n_23378;
assign n_23380 =  x_2687 & ~n_23379;
assign n_23381 = ~x_2687 &  n_23379;
assign n_23382 = ~n_23380 & ~n_23381;
assign n_23383 =  x_2686 & ~n_23310;
assign n_23384 =  i_20 &  n_23310;
assign n_23385 = ~n_23383 & ~n_23384;
assign n_23386 =  x_2686 & ~n_23385;
assign n_23387 = ~x_2686 &  n_23385;
assign n_23388 = ~n_23386 & ~n_23387;
assign n_23389 =  x_2685 & ~n_23310;
assign n_23390 =  i_19 &  n_23310;
assign n_23391 = ~n_23389 & ~n_23390;
assign n_23392 =  x_2685 & ~n_23391;
assign n_23393 = ~x_2685 &  n_23391;
assign n_23394 = ~n_23392 & ~n_23393;
assign n_23395 =  x_2684 & ~n_23310;
assign n_23396 =  i_18 &  n_23310;
assign n_23397 = ~n_23395 & ~n_23396;
assign n_23398 =  x_2684 & ~n_23397;
assign n_23399 = ~x_2684 &  n_23397;
assign n_23400 = ~n_23398 & ~n_23399;
assign n_23401 =  x_2683 & ~n_23310;
assign n_23402 =  i_17 &  n_23310;
assign n_23403 = ~n_23401 & ~n_23402;
assign n_23404 =  x_2683 & ~n_23403;
assign n_23405 = ~x_2683 &  n_23403;
assign n_23406 = ~n_23404 & ~n_23405;
assign n_23407 =  x_2682 & ~n_23310;
assign n_23408 =  i_16 &  n_23310;
assign n_23409 = ~n_23407 & ~n_23408;
assign n_23410 =  x_2682 & ~n_23409;
assign n_23411 = ~x_2682 &  n_23409;
assign n_23412 = ~n_23410 & ~n_23411;
assign n_23413 =  x_2681 & ~n_23310;
assign n_23414 =  i_15 &  n_23310;
assign n_23415 = ~n_23413 & ~n_23414;
assign n_23416 =  x_2681 & ~n_23415;
assign n_23417 = ~x_2681 &  n_23415;
assign n_23418 = ~n_23416 & ~n_23417;
assign n_23419 =  x_2680 & ~n_23310;
assign n_23420 =  i_14 &  n_23310;
assign n_23421 = ~n_23419 & ~n_23420;
assign n_23422 =  x_2680 & ~n_23421;
assign n_23423 = ~x_2680 &  n_23421;
assign n_23424 = ~n_23422 & ~n_23423;
assign n_23425 =  x_2679 & ~n_23310;
assign n_23426 =  i_13 &  n_23310;
assign n_23427 = ~n_23425 & ~n_23426;
assign n_23428 =  x_2679 & ~n_23427;
assign n_23429 = ~x_2679 &  n_23427;
assign n_23430 = ~n_23428 & ~n_23429;
assign n_23431 =  x_2678 & ~n_23310;
assign n_23432 =  i_12 &  n_23310;
assign n_23433 = ~n_23431 & ~n_23432;
assign n_23434 =  x_2678 & ~n_23433;
assign n_23435 = ~x_2678 &  n_23433;
assign n_23436 = ~n_23434 & ~n_23435;
assign n_23437 =  x_2677 & ~n_23310;
assign n_23438 =  i_11 &  n_23310;
assign n_23439 = ~n_23437 & ~n_23438;
assign n_23440 =  x_2677 & ~n_23439;
assign n_23441 = ~x_2677 &  n_23439;
assign n_23442 = ~n_23440 & ~n_23441;
assign n_23443 =  x_2676 & ~n_23310;
assign n_23444 =  i_10 &  n_23310;
assign n_23445 = ~n_23443 & ~n_23444;
assign n_23446 =  x_2676 & ~n_23445;
assign n_23447 = ~x_2676 &  n_23445;
assign n_23448 = ~n_23446 & ~n_23447;
assign n_23449 =  x_2675 & ~n_23310;
assign n_23450 =  i_9 &  n_23310;
assign n_23451 = ~n_23449 & ~n_23450;
assign n_23452 =  x_2675 & ~n_23451;
assign n_23453 = ~x_2675 &  n_23451;
assign n_23454 = ~n_23452 & ~n_23453;
assign n_23455 =  x_2674 & ~n_23310;
assign n_23456 =  i_8 &  n_23310;
assign n_23457 = ~n_23455 & ~n_23456;
assign n_23458 =  x_2674 & ~n_23457;
assign n_23459 = ~x_2674 &  n_23457;
assign n_23460 = ~n_23458 & ~n_23459;
assign n_23461 =  x_2673 & ~n_23310;
assign n_23462 =  i_7 &  n_23310;
assign n_23463 = ~n_23461 & ~n_23462;
assign n_23464 =  x_2673 & ~n_23463;
assign n_23465 = ~x_2673 &  n_23463;
assign n_23466 = ~n_23464 & ~n_23465;
assign n_23467 =  x_2672 & ~n_23310;
assign n_23468 =  i_6 &  n_23310;
assign n_23469 = ~n_23467 & ~n_23468;
assign n_23470 =  x_2672 & ~n_23469;
assign n_23471 = ~x_2672 &  n_23469;
assign n_23472 = ~n_23470 & ~n_23471;
assign n_23473 =  x_2671 & ~n_23310;
assign n_23474 =  i_5 &  n_23310;
assign n_23475 = ~n_23473 & ~n_23474;
assign n_23476 =  x_2671 & ~n_23475;
assign n_23477 = ~x_2671 &  n_23475;
assign n_23478 = ~n_23476 & ~n_23477;
assign n_23479 =  x_2670 & ~n_23310;
assign n_23480 =  i_4 &  n_23310;
assign n_23481 = ~n_23479 & ~n_23480;
assign n_23482 =  x_2670 & ~n_23481;
assign n_23483 = ~x_2670 &  n_23481;
assign n_23484 = ~n_23482 & ~n_23483;
assign n_23485 =  x_2669 & ~n_23310;
assign n_23486 =  i_3 &  n_23310;
assign n_23487 = ~n_23485 & ~n_23486;
assign n_23488 =  x_2669 & ~n_23487;
assign n_23489 = ~x_2669 &  n_23487;
assign n_23490 = ~n_23488 & ~n_23489;
assign n_23491 =  x_2668 & ~n_23310;
assign n_23492 =  i_2 &  n_23310;
assign n_23493 = ~n_23491 & ~n_23492;
assign n_23494 =  x_2668 & ~n_23493;
assign n_23495 = ~x_2668 &  n_23493;
assign n_23496 = ~n_23494 & ~n_23495;
assign n_23497 =  x_2667 & ~n_23310;
assign n_23498 =  i_1 &  n_23310;
assign n_23499 = ~n_23497 & ~n_23498;
assign n_23500 =  x_2667 & ~n_23499;
assign n_23501 = ~x_2667 &  n_23499;
assign n_23502 = ~n_23500 & ~n_23501;
assign n_23503 =  n_3858 &  n_8;
assign n_23504 =  x_39 &  n_23503;
assign n_23505 =  x_2666 & ~n_23504;
assign n_23506 =  i_32 &  n_23504;
assign n_23507 = ~n_23505 & ~n_23506;
assign n_23508 =  x_2666 & ~n_23507;
assign n_23509 = ~x_2666 &  n_23507;
assign n_23510 = ~n_23508 & ~n_23509;
assign n_23511 =  x_2665 & ~n_23504;
assign n_23512 =  i_31 &  n_23504;
assign n_23513 = ~n_23511 & ~n_23512;
assign n_23514 =  x_2665 & ~n_23513;
assign n_23515 = ~x_2665 &  n_23513;
assign n_23516 = ~n_23514 & ~n_23515;
assign n_23517 =  x_2664 & ~n_23504;
assign n_23518 =  i_30 &  n_23504;
assign n_23519 = ~n_23517 & ~n_23518;
assign n_23520 =  x_2664 & ~n_23519;
assign n_23521 = ~x_2664 &  n_23519;
assign n_23522 = ~n_23520 & ~n_23521;
assign n_23523 =  x_2663 & ~n_23504;
assign n_23524 =  i_29 &  n_23504;
assign n_23525 = ~n_23523 & ~n_23524;
assign n_23526 =  x_2663 & ~n_23525;
assign n_23527 = ~x_2663 &  n_23525;
assign n_23528 = ~n_23526 & ~n_23527;
assign n_23529 =  x_2662 & ~n_23504;
assign n_23530 =  i_28 &  n_23504;
assign n_23531 = ~n_23529 & ~n_23530;
assign n_23532 =  x_2662 & ~n_23531;
assign n_23533 = ~x_2662 &  n_23531;
assign n_23534 = ~n_23532 & ~n_23533;
assign n_23535 =  x_2661 & ~n_23504;
assign n_23536 =  i_27 &  n_23504;
assign n_23537 = ~n_23535 & ~n_23536;
assign n_23538 =  x_2661 & ~n_23537;
assign n_23539 = ~x_2661 &  n_23537;
assign n_23540 = ~n_23538 & ~n_23539;
assign n_23541 =  x_2660 & ~n_23504;
assign n_23542 =  i_26 &  n_23504;
assign n_23543 = ~n_23541 & ~n_23542;
assign n_23544 =  x_2660 & ~n_23543;
assign n_23545 = ~x_2660 &  n_23543;
assign n_23546 = ~n_23544 & ~n_23545;
assign n_23547 =  x_2659 & ~n_23504;
assign n_23548 =  i_25 &  n_23504;
assign n_23549 = ~n_23547 & ~n_23548;
assign n_23550 =  x_2659 & ~n_23549;
assign n_23551 = ~x_2659 &  n_23549;
assign n_23552 = ~n_23550 & ~n_23551;
assign n_23553 =  x_2658 & ~n_23504;
assign n_23554 =  i_24 &  n_23504;
assign n_23555 = ~n_23553 & ~n_23554;
assign n_23556 =  x_2658 & ~n_23555;
assign n_23557 = ~x_2658 &  n_23555;
assign n_23558 = ~n_23556 & ~n_23557;
assign n_23559 =  x_2657 & ~n_23504;
assign n_23560 =  i_23 &  n_23504;
assign n_23561 = ~n_23559 & ~n_23560;
assign n_23562 =  x_2657 & ~n_23561;
assign n_23563 = ~x_2657 &  n_23561;
assign n_23564 = ~n_23562 & ~n_23563;
assign n_23565 =  x_2656 & ~n_23504;
assign n_23566 =  i_22 &  n_23504;
assign n_23567 = ~n_23565 & ~n_23566;
assign n_23568 =  x_2656 & ~n_23567;
assign n_23569 = ~x_2656 &  n_23567;
assign n_23570 = ~n_23568 & ~n_23569;
assign n_23571 =  x_2655 & ~n_23504;
assign n_23572 =  i_21 &  n_23504;
assign n_23573 = ~n_23571 & ~n_23572;
assign n_23574 =  x_2655 & ~n_23573;
assign n_23575 = ~x_2655 &  n_23573;
assign n_23576 = ~n_23574 & ~n_23575;
assign n_23577 =  x_2654 & ~n_23504;
assign n_23578 =  i_20 &  n_23504;
assign n_23579 = ~n_23577 & ~n_23578;
assign n_23580 =  x_2654 & ~n_23579;
assign n_23581 = ~x_2654 &  n_23579;
assign n_23582 = ~n_23580 & ~n_23581;
assign n_23583 =  x_2653 & ~n_23504;
assign n_23584 =  i_19 &  n_23504;
assign n_23585 = ~n_23583 & ~n_23584;
assign n_23586 =  x_2653 & ~n_23585;
assign n_23587 = ~x_2653 &  n_23585;
assign n_23588 = ~n_23586 & ~n_23587;
assign n_23589 =  x_2652 & ~n_23504;
assign n_23590 =  i_18 &  n_23504;
assign n_23591 = ~n_23589 & ~n_23590;
assign n_23592 =  x_2652 & ~n_23591;
assign n_23593 = ~x_2652 &  n_23591;
assign n_23594 = ~n_23592 & ~n_23593;
assign n_23595 =  x_2651 & ~n_23504;
assign n_23596 =  i_17 &  n_23504;
assign n_23597 = ~n_23595 & ~n_23596;
assign n_23598 =  x_2651 & ~n_23597;
assign n_23599 = ~x_2651 &  n_23597;
assign n_23600 = ~n_23598 & ~n_23599;
assign n_23601 =  x_2650 & ~n_23504;
assign n_23602 =  i_16 &  n_23504;
assign n_23603 = ~n_23601 & ~n_23602;
assign n_23604 =  x_2650 & ~n_23603;
assign n_23605 = ~x_2650 &  n_23603;
assign n_23606 = ~n_23604 & ~n_23605;
assign n_23607 =  x_2649 & ~n_23504;
assign n_23608 =  i_15 &  n_23504;
assign n_23609 = ~n_23607 & ~n_23608;
assign n_23610 =  x_2649 & ~n_23609;
assign n_23611 = ~x_2649 &  n_23609;
assign n_23612 = ~n_23610 & ~n_23611;
assign n_23613 =  x_2648 & ~n_23504;
assign n_23614 =  i_14 &  n_23504;
assign n_23615 = ~n_23613 & ~n_23614;
assign n_23616 =  x_2648 & ~n_23615;
assign n_23617 = ~x_2648 &  n_23615;
assign n_23618 = ~n_23616 & ~n_23617;
assign n_23619 =  x_2647 & ~n_23504;
assign n_23620 =  i_13 &  n_23504;
assign n_23621 = ~n_23619 & ~n_23620;
assign n_23622 =  x_2647 & ~n_23621;
assign n_23623 = ~x_2647 &  n_23621;
assign n_23624 = ~n_23622 & ~n_23623;
assign n_23625 =  x_2646 & ~n_23504;
assign n_23626 =  i_12 &  n_23504;
assign n_23627 = ~n_23625 & ~n_23626;
assign n_23628 =  x_2646 & ~n_23627;
assign n_23629 = ~x_2646 &  n_23627;
assign n_23630 = ~n_23628 & ~n_23629;
assign n_23631 =  x_2645 & ~n_23504;
assign n_23632 =  i_11 &  n_23504;
assign n_23633 = ~n_23631 & ~n_23632;
assign n_23634 =  x_2645 & ~n_23633;
assign n_23635 = ~x_2645 &  n_23633;
assign n_23636 = ~n_23634 & ~n_23635;
assign n_23637 =  x_2644 & ~n_23504;
assign n_23638 =  i_10 &  n_23504;
assign n_23639 = ~n_23637 & ~n_23638;
assign n_23640 =  x_2644 & ~n_23639;
assign n_23641 = ~x_2644 &  n_23639;
assign n_23642 = ~n_23640 & ~n_23641;
assign n_23643 =  x_2643 & ~n_23504;
assign n_23644 =  i_9 &  n_23504;
assign n_23645 = ~n_23643 & ~n_23644;
assign n_23646 =  x_2643 & ~n_23645;
assign n_23647 = ~x_2643 &  n_23645;
assign n_23648 = ~n_23646 & ~n_23647;
assign n_23649 =  x_2642 & ~n_23504;
assign n_23650 =  i_8 &  n_23504;
assign n_23651 = ~n_23649 & ~n_23650;
assign n_23652 =  x_2642 & ~n_23651;
assign n_23653 = ~x_2642 &  n_23651;
assign n_23654 = ~n_23652 & ~n_23653;
assign n_23655 =  x_2641 & ~n_23504;
assign n_23656 =  i_7 &  n_23504;
assign n_23657 = ~n_23655 & ~n_23656;
assign n_23658 =  x_2641 & ~n_23657;
assign n_23659 = ~x_2641 &  n_23657;
assign n_23660 = ~n_23658 & ~n_23659;
assign n_23661 =  x_2640 & ~n_23504;
assign n_23662 =  i_6 &  n_23504;
assign n_23663 = ~n_23661 & ~n_23662;
assign n_23664 =  x_2640 & ~n_23663;
assign n_23665 = ~x_2640 &  n_23663;
assign n_23666 = ~n_23664 & ~n_23665;
assign n_23667 =  x_2639 & ~n_23504;
assign n_23668 =  i_5 &  n_23504;
assign n_23669 = ~n_23667 & ~n_23668;
assign n_23670 =  x_2639 & ~n_23669;
assign n_23671 = ~x_2639 &  n_23669;
assign n_23672 = ~n_23670 & ~n_23671;
assign n_23673 =  x_2638 & ~n_23504;
assign n_23674 =  i_4 &  n_23504;
assign n_23675 = ~n_23673 & ~n_23674;
assign n_23676 =  x_2638 & ~n_23675;
assign n_23677 = ~x_2638 &  n_23675;
assign n_23678 = ~n_23676 & ~n_23677;
assign n_23679 =  x_2637 & ~n_23504;
assign n_23680 =  i_3 &  n_23504;
assign n_23681 = ~n_23679 & ~n_23680;
assign n_23682 =  x_2637 & ~n_23681;
assign n_23683 = ~x_2637 &  n_23681;
assign n_23684 = ~n_23682 & ~n_23683;
assign n_23685 =  x_2636 & ~n_23504;
assign n_23686 =  i_2 &  n_23504;
assign n_23687 = ~n_23685 & ~n_23686;
assign n_23688 =  x_2636 & ~n_23687;
assign n_23689 = ~x_2636 &  n_23687;
assign n_23690 = ~n_23688 & ~n_23689;
assign n_23691 =  x_2635 & ~n_23504;
assign n_23692 =  i_1 &  n_23504;
assign n_23693 = ~n_23691 & ~n_23692;
assign n_23694 =  x_2635 & ~n_23693;
assign n_23695 = ~x_2635 &  n_23693;
assign n_23696 = ~n_23694 & ~n_23695;
assign n_23697 =  n_4 &  n_587;
assign n_23698 =  n_1903 &  n_23697;
assign n_23699 =  x_2634 & ~n_23698;
assign n_23700 =  i_32 &  n_23698;
assign n_23701 = ~n_23699 & ~n_23700;
assign n_23702 =  x_2634 & ~n_23701;
assign n_23703 = ~x_2634 &  n_23701;
assign n_23704 = ~n_23702 & ~n_23703;
assign n_23705 =  x_2633 & ~n_23698;
assign n_23706 =  i_31 &  n_23698;
assign n_23707 = ~n_23705 & ~n_23706;
assign n_23708 =  x_2633 & ~n_23707;
assign n_23709 = ~x_2633 &  n_23707;
assign n_23710 = ~n_23708 & ~n_23709;
assign n_23711 =  x_2632 & ~n_23698;
assign n_23712 =  i_30 &  n_23698;
assign n_23713 = ~n_23711 & ~n_23712;
assign n_23714 =  x_2632 & ~n_23713;
assign n_23715 = ~x_2632 &  n_23713;
assign n_23716 = ~n_23714 & ~n_23715;
assign n_23717 =  x_2631 & ~n_23698;
assign n_23718 =  i_29 &  n_23698;
assign n_23719 = ~n_23717 & ~n_23718;
assign n_23720 =  x_2631 & ~n_23719;
assign n_23721 = ~x_2631 &  n_23719;
assign n_23722 = ~n_23720 & ~n_23721;
assign n_23723 =  x_2630 & ~n_23698;
assign n_23724 =  i_28 &  n_23698;
assign n_23725 = ~n_23723 & ~n_23724;
assign n_23726 =  x_2630 & ~n_23725;
assign n_23727 = ~x_2630 &  n_23725;
assign n_23728 = ~n_23726 & ~n_23727;
assign n_23729 =  x_2629 & ~n_23698;
assign n_23730 =  i_27 &  n_23698;
assign n_23731 = ~n_23729 & ~n_23730;
assign n_23732 =  x_2629 & ~n_23731;
assign n_23733 = ~x_2629 &  n_23731;
assign n_23734 = ~n_23732 & ~n_23733;
assign n_23735 =  x_2628 & ~n_23698;
assign n_23736 =  i_26 &  n_23698;
assign n_23737 = ~n_23735 & ~n_23736;
assign n_23738 =  x_2628 & ~n_23737;
assign n_23739 = ~x_2628 &  n_23737;
assign n_23740 = ~n_23738 & ~n_23739;
assign n_23741 =  x_2627 & ~n_23698;
assign n_23742 =  i_25 &  n_23698;
assign n_23743 = ~n_23741 & ~n_23742;
assign n_23744 =  x_2627 & ~n_23743;
assign n_23745 = ~x_2627 &  n_23743;
assign n_23746 = ~n_23744 & ~n_23745;
assign n_23747 =  x_2626 & ~n_23698;
assign n_23748 =  i_24 &  n_23698;
assign n_23749 = ~n_23747 & ~n_23748;
assign n_23750 =  x_2626 & ~n_23749;
assign n_23751 = ~x_2626 &  n_23749;
assign n_23752 = ~n_23750 & ~n_23751;
assign n_23753 =  x_2625 & ~n_23698;
assign n_23754 =  i_23 &  n_23698;
assign n_23755 = ~n_23753 & ~n_23754;
assign n_23756 =  x_2625 & ~n_23755;
assign n_23757 = ~x_2625 &  n_23755;
assign n_23758 = ~n_23756 & ~n_23757;
assign n_23759 =  x_2624 & ~n_23698;
assign n_23760 =  i_22 &  n_23698;
assign n_23761 = ~n_23759 & ~n_23760;
assign n_23762 =  x_2624 & ~n_23761;
assign n_23763 = ~x_2624 &  n_23761;
assign n_23764 = ~n_23762 & ~n_23763;
assign n_23765 =  x_2623 & ~n_23698;
assign n_23766 =  i_21 &  n_23698;
assign n_23767 = ~n_23765 & ~n_23766;
assign n_23768 =  x_2623 & ~n_23767;
assign n_23769 = ~x_2623 &  n_23767;
assign n_23770 = ~n_23768 & ~n_23769;
assign n_23771 =  x_2622 & ~n_23698;
assign n_23772 =  i_20 &  n_23698;
assign n_23773 = ~n_23771 & ~n_23772;
assign n_23774 =  x_2622 & ~n_23773;
assign n_23775 = ~x_2622 &  n_23773;
assign n_23776 = ~n_23774 & ~n_23775;
assign n_23777 =  x_2621 & ~n_23698;
assign n_23778 =  i_19 &  n_23698;
assign n_23779 = ~n_23777 & ~n_23778;
assign n_23780 =  x_2621 & ~n_23779;
assign n_23781 = ~x_2621 &  n_23779;
assign n_23782 = ~n_23780 & ~n_23781;
assign n_23783 =  x_2620 & ~n_23698;
assign n_23784 =  i_18 &  n_23698;
assign n_23785 = ~n_23783 & ~n_23784;
assign n_23786 =  x_2620 & ~n_23785;
assign n_23787 = ~x_2620 &  n_23785;
assign n_23788 = ~n_23786 & ~n_23787;
assign n_23789 =  x_2619 & ~n_23698;
assign n_23790 =  i_17 &  n_23698;
assign n_23791 = ~n_23789 & ~n_23790;
assign n_23792 =  x_2619 & ~n_23791;
assign n_23793 = ~x_2619 &  n_23791;
assign n_23794 = ~n_23792 & ~n_23793;
assign n_23795 =  x_2618 & ~n_23698;
assign n_23796 =  i_16 &  n_23698;
assign n_23797 = ~n_23795 & ~n_23796;
assign n_23798 =  x_2618 & ~n_23797;
assign n_23799 = ~x_2618 &  n_23797;
assign n_23800 = ~n_23798 & ~n_23799;
assign n_23801 =  x_2617 & ~n_23698;
assign n_23802 =  i_15 &  n_23698;
assign n_23803 = ~n_23801 & ~n_23802;
assign n_23804 =  x_2617 & ~n_23803;
assign n_23805 = ~x_2617 &  n_23803;
assign n_23806 = ~n_23804 & ~n_23805;
assign n_23807 =  x_2616 & ~n_23698;
assign n_23808 =  i_14 &  n_23698;
assign n_23809 = ~n_23807 & ~n_23808;
assign n_23810 =  x_2616 & ~n_23809;
assign n_23811 = ~x_2616 &  n_23809;
assign n_23812 = ~n_23810 & ~n_23811;
assign n_23813 =  x_2615 & ~n_23698;
assign n_23814 =  i_13 &  n_23698;
assign n_23815 = ~n_23813 & ~n_23814;
assign n_23816 =  x_2615 & ~n_23815;
assign n_23817 = ~x_2615 &  n_23815;
assign n_23818 = ~n_23816 & ~n_23817;
assign n_23819 =  x_2614 & ~n_23698;
assign n_23820 =  i_12 &  n_23698;
assign n_23821 = ~n_23819 & ~n_23820;
assign n_23822 =  x_2614 & ~n_23821;
assign n_23823 = ~x_2614 &  n_23821;
assign n_23824 = ~n_23822 & ~n_23823;
assign n_23825 =  x_2613 & ~n_23698;
assign n_23826 =  i_11 &  n_23698;
assign n_23827 = ~n_23825 & ~n_23826;
assign n_23828 =  x_2613 & ~n_23827;
assign n_23829 = ~x_2613 &  n_23827;
assign n_23830 = ~n_23828 & ~n_23829;
assign n_23831 =  x_2612 & ~n_23698;
assign n_23832 =  i_10 &  n_23698;
assign n_23833 = ~n_23831 & ~n_23832;
assign n_23834 =  x_2612 & ~n_23833;
assign n_23835 = ~x_2612 &  n_23833;
assign n_23836 = ~n_23834 & ~n_23835;
assign n_23837 =  x_2611 & ~n_23698;
assign n_23838 =  i_9 &  n_23698;
assign n_23839 = ~n_23837 & ~n_23838;
assign n_23840 =  x_2611 & ~n_23839;
assign n_23841 = ~x_2611 &  n_23839;
assign n_23842 = ~n_23840 & ~n_23841;
assign n_23843 =  x_2610 & ~n_23698;
assign n_23844 =  i_8 &  n_23698;
assign n_23845 = ~n_23843 & ~n_23844;
assign n_23846 =  x_2610 & ~n_23845;
assign n_23847 = ~x_2610 &  n_23845;
assign n_23848 = ~n_23846 & ~n_23847;
assign n_23849 =  x_2609 & ~n_23698;
assign n_23850 =  i_7 &  n_23698;
assign n_23851 = ~n_23849 & ~n_23850;
assign n_23852 =  x_2609 & ~n_23851;
assign n_23853 = ~x_2609 &  n_23851;
assign n_23854 = ~n_23852 & ~n_23853;
assign n_23855 =  x_2608 & ~n_23698;
assign n_23856 =  i_6 &  n_23698;
assign n_23857 = ~n_23855 & ~n_23856;
assign n_23858 =  x_2608 & ~n_23857;
assign n_23859 = ~x_2608 &  n_23857;
assign n_23860 = ~n_23858 & ~n_23859;
assign n_23861 =  x_2607 & ~n_23698;
assign n_23862 =  i_5 &  n_23698;
assign n_23863 = ~n_23861 & ~n_23862;
assign n_23864 =  x_2607 & ~n_23863;
assign n_23865 = ~x_2607 &  n_23863;
assign n_23866 = ~n_23864 & ~n_23865;
assign n_23867 =  x_2606 & ~n_23698;
assign n_23868 =  i_4 &  n_23698;
assign n_23869 = ~n_23867 & ~n_23868;
assign n_23870 =  x_2606 & ~n_23869;
assign n_23871 = ~x_2606 &  n_23869;
assign n_23872 = ~n_23870 & ~n_23871;
assign n_23873 =  x_2605 & ~n_23698;
assign n_23874 =  i_3 &  n_23698;
assign n_23875 = ~n_23873 & ~n_23874;
assign n_23876 =  x_2605 & ~n_23875;
assign n_23877 = ~x_2605 &  n_23875;
assign n_23878 = ~n_23876 & ~n_23877;
assign n_23879 =  x_2604 & ~n_23698;
assign n_23880 =  i_2 &  n_23698;
assign n_23881 = ~n_23879 & ~n_23880;
assign n_23882 =  x_2604 & ~n_23881;
assign n_23883 = ~x_2604 &  n_23881;
assign n_23884 = ~n_23882 & ~n_23883;
assign n_23885 =  x_2603 & ~n_23698;
assign n_23886 =  i_1 &  n_23698;
assign n_23887 = ~n_23885 & ~n_23886;
assign n_23888 =  x_2603 & ~n_23887;
assign n_23889 = ~x_2603 &  n_23887;
assign n_23890 = ~n_23888 & ~n_23889;
assign n_23891 =  n_389 &  n_982;
assign n_23892 = ~x_39 &  n_23891;
assign n_23893 =  n_2301 &  n_23892;
assign n_23894 =  n_3663 &  n_23891;
assign n_23895 = ~n_23893 & ~n_23894;
assign n_23896 =  x_2602 &  n_23895;
assign n_23897 = ~n_3664 & ~n_12420;
assign n_23898 = ~n_23897 &  n_23891;
assign n_23899 = ~n_23896 & ~n_23898;
assign n_23900 =  x_2602 & ~n_23899;
assign n_23901 = ~x_2602 &  n_23899;
assign n_23902 = ~n_23900 & ~n_23901;
assign n_23903 =  x_2601 &  n_23895;
assign n_23904 =  x_2601 &  n_23903;
assign n_23905 = ~x_2601 & ~n_23903;
assign n_23906 = ~n_23904 & ~n_23905;
assign n_23907 =  x_2600 &  n_23895;
assign n_23908 =  x_2600 &  n_23907;
assign n_23909 = ~x_2600 & ~n_23907;
assign n_23910 = ~n_23908 & ~n_23909;
assign n_23911 =  x_2599 &  n_23895;
assign n_23912 =  x_2599 &  n_23911;
assign n_23913 = ~x_2599 & ~n_23911;
assign n_23914 = ~n_23912 & ~n_23913;
assign n_23915 =  x_2598 &  n_23895;
assign n_23916 =  x_2598 &  n_23915;
assign n_23917 = ~x_2598 & ~n_23915;
assign n_23918 = ~n_23916 & ~n_23917;
assign n_23919 =  x_2597 &  n_23895;
assign n_23920 =  x_2597 &  n_23919;
assign n_23921 = ~x_2597 & ~n_23919;
assign n_23922 = ~n_23920 & ~n_23921;
assign n_23923 =  x_2596 &  n_23895;
assign n_23924 =  x_2596 &  n_23923;
assign n_23925 = ~x_2596 & ~n_23923;
assign n_23926 = ~n_23924 & ~n_23925;
assign n_23927 =  x_2595 &  n_23895;
assign n_23928 =  x_2595 &  n_23927;
assign n_23929 = ~x_2595 & ~n_23927;
assign n_23930 = ~n_23928 & ~n_23929;
assign n_23931 =  x_2594 &  n_23895;
assign n_23932 =  x_2594 &  n_23931;
assign n_23933 = ~x_2594 & ~n_23931;
assign n_23934 = ~n_23932 & ~n_23933;
assign n_23935 =  x_2593 &  n_23895;
assign n_23936 =  x_2593 &  n_23935;
assign n_23937 = ~x_2593 & ~n_23935;
assign n_23938 = ~n_23936 & ~n_23937;
assign n_23939 =  x_2592 &  n_23895;
assign n_23940 =  x_2592 &  n_23939;
assign n_23941 = ~x_2592 & ~n_23939;
assign n_23942 = ~n_23940 & ~n_23941;
assign n_23943 =  x_2591 &  n_23895;
assign n_23944 =  x_2591 &  n_23943;
assign n_23945 = ~x_2591 & ~n_23943;
assign n_23946 = ~n_23944 & ~n_23945;
assign n_23947 =  x_2590 &  n_23895;
assign n_23948 =  x_2590 &  n_23947;
assign n_23949 = ~x_2590 & ~n_23947;
assign n_23950 = ~n_23948 & ~n_23949;
assign n_23951 =  x_2589 &  n_23895;
assign n_23952 =  x_2589 &  n_23951;
assign n_23953 = ~x_2589 & ~n_23951;
assign n_23954 = ~n_23952 & ~n_23953;
assign n_23955 =  x_2588 &  n_23895;
assign n_23956 =  x_2588 &  n_23955;
assign n_23957 = ~x_2588 & ~n_23955;
assign n_23958 = ~n_23956 & ~n_23957;
assign n_23959 =  x_2587 &  n_23895;
assign n_23960 =  x_2587 &  n_23959;
assign n_23961 = ~x_2587 & ~n_23959;
assign n_23962 = ~n_23960 & ~n_23961;
assign n_23963 =  x_2586 &  n_23895;
assign n_23964 =  x_2586 &  n_23963;
assign n_23965 = ~x_2586 & ~n_23963;
assign n_23966 = ~n_23964 & ~n_23965;
assign n_23967 =  x_2585 &  n_23895;
assign n_23968 =  x_2585 &  n_23967;
assign n_23969 = ~x_2585 & ~n_23967;
assign n_23970 = ~n_23968 & ~n_23969;
assign n_23971 =  x_2584 &  n_23895;
assign n_23972 =  x_2584 &  n_23971;
assign n_23973 = ~x_2584 & ~n_23971;
assign n_23974 = ~n_23972 & ~n_23973;
assign n_23975 =  x_2583 &  n_23895;
assign n_23976 =  x_2583 &  n_23975;
assign n_23977 = ~x_2583 & ~n_23975;
assign n_23978 = ~n_23976 & ~n_23977;
assign n_23979 =  x_2582 &  n_23895;
assign n_23980 =  x_2582 &  n_23979;
assign n_23981 = ~x_2582 & ~n_23979;
assign n_23982 = ~n_23980 & ~n_23981;
assign n_23983 =  x_2581 &  n_23895;
assign n_23984 =  x_2581 &  n_23983;
assign n_23985 = ~x_2581 & ~n_23983;
assign n_23986 = ~n_23984 & ~n_23985;
assign n_23987 =  x_2580 &  n_23895;
assign n_23988 =  x_2580 &  n_23987;
assign n_23989 = ~x_2580 & ~n_23987;
assign n_23990 = ~n_23988 & ~n_23989;
assign n_23991 =  x_2579 &  n_23895;
assign n_23992 =  x_2579 &  n_23991;
assign n_23993 = ~x_2579 & ~n_23991;
assign n_23994 = ~n_23992 & ~n_23993;
assign n_23995 =  x_2578 &  n_23895;
assign n_23996 =  x_2578 &  n_23995;
assign n_23997 = ~x_2578 & ~n_23995;
assign n_23998 = ~n_23996 & ~n_23997;
assign n_23999 =  x_2577 &  n_23895;
assign n_24000 =  x_2577 &  n_23999;
assign n_24001 = ~x_2577 & ~n_23999;
assign n_24002 = ~n_24000 & ~n_24001;
assign n_24003 =  x_2576 &  n_23895;
assign n_24004 =  x_2576 &  n_24003;
assign n_24005 = ~x_2576 & ~n_24003;
assign n_24006 = ~n_24004 & ~n_24005;
assign n_24007 =  x_2575 &  n_23895;
assign n_24008 =  x_2575 &  n_24007;
assign n_24009 = ~x_2575 & ~n_24007;
assign n_24010 = ~n_24008 & ~n_24009;
assign n_24011 =  x_2574 &  n_23895;
assign n_24012 =  x_2574 &  n_24011;
assign n_24013 = ~x_2574 & ~n_24011;
assign n_24014 = ~n_24012 & ~n_24013;
assign n_24015 =  x_2573 &  n_23895;
assign n_24016 =  x_2573 &  n_24015;
assign n_24017 = ~x_2573 & ~n_24015;
assign n_24018 = ~n_24016 & ~n_24017;
assign n_24019 =  x_2572 &  n_23895;
assign n_24020 =  x_2572 &  n_24019;
assign n_24021 = ~x_2572 & ~n_24019;
assign n_24022 = ~n_24020 & ~n_24021;
assign n_24023 =  x_2571 &  n_23895;
assign n_24024 =  x_2571 &  n_24023;
assign n_24025 = ~x_2571 & ~n_24023;
assign n_24026 = ~n_24024 & ~n_24025;
assign n_24027 =  n_3469 &  n_2499;
assign n_24028 =  x_2570 & ~n_24027;
assign n_24029 =  i_32 &  n_24027;
assign n_24030 = ~n_24028 & ~n_24029;
assign n_24031 =  x_2570 & ~n_24030;
assign n_24032 = ~x_2570 &  n_24030;
assign n_24033 = ~n_24031 & ~n_24032;
assign n_24034 =  x_2569 & ~n_24027;
assign n_24035 =  i_31 &  n_24027;
assign n_24036 = ~n_24034 & ~n_24035;
assign n_24037 =  x_2569 & ~n_24036;
assign n_24038 = ~x_2569 &  n_24036;
assign n_24039 = ~n_24037 & ~n_24038;
assign n_24040 =  x_2568 & ~n_24027;
assign n_24041 =  i_30 &  n_24027;
assign n_24042 = ~n_24040 & ~n_24041;
assign n_24043 =  x_2568 & ~n_24042;
assign n_24044 = ~x_2568 &  n_24042;
assign n_24045 = ~n_24043 & ~n_24044;
assign n_24046 =  x_2567 & ~n_24027;
assign n_24047 =  i_29 &  n_24027;
assign n_24048 = ~n_24046 & ~n_24047;
assign n_24049 =  x_2567 & ~n_24048;
assign n_24050 = ~x_2567 &  n_24048;
assign n_24051 = ~n_24049 & ~n_24050;
assign n_24052 =  x_2566 & ~n_24027;
assign n_24053 =  i_28 &  n_24027;
assign n_24054 = ~n_24052 & ~n_24053;
assign n_24055 =  x_2566 & ~n_24054;
assign n_24056 = ~x_2566 &  n_24054;
assign n_24057 = ~n_24055 & ~n_24056;
assign n_24058 =  x_2565 & ~n_24027;
assign n_24059 =  i_27 &  n_24027;
assign n_24060 = ~n_24058 & ~n_24059;
assign n_24061 =  x_2565 & ~n_24060;
assign n_24062 = ~x_2565 &  n_24060;
assign n_24063 = ~n_24061 & ~n_24062;
assign n_24064 =  x_2564 & ~n_24027;
assign n_24065 =  i_26 &  n_24027;
assign n_24066 = ~n_24064 & ~n_24065;
assign n_24067 =  x_2564 & ~n_24066;
assign n_24068 = ~x_2564 &  n_24066;
assign n_24069 = ~n_24067 & ~n_24068;
assign n_24070 =  x_2563 & ~n_24027;
assign n_24071 =  i_25 &  n_24027;
assign n_24072 = ~n_24070 & ~n_24071;
assign n_24073 =  x_2563 & ~n_24072;
assign n_24074 = ~x_2563 &  n_24072;
assign n_24075 = ~n_24073 & ~n_24074;
assign n_24076 =  x_2562 & ~n_24027;
assign n_24077 =  i_24 &  n_24027;
assign n_24078 = ~n_24076 & ~n_24077;
assign n_24079 =  x_2562 & ~n_24078;
assign n_24080 = ~x_2562 &  n_24078;
assign n_24081 = ~n_24079 & ~n_24080;
assign n_24082 =  x_2561 & ~n_24027;
assign n_24083 =  i_23 &  n_24027;
assign n_24084 = ~n_24082 & ~n_24083;
assign n_24085 =  x_2561 & ~n_24084;
assign n_24086 = ~x_2561 &  n_24084;
assign n_24087 = ~n_24085 & ~n_24086;
assign n_24088 =  x_2560 & ~n_24027;
assign n_24089 =  i_22 &  n_24027;
assign n_24090 = ~n_24088 & ~n_24089;
assign n_24091 =  x_2560 & ~n_24090;
assign n_24092 = ~x_2560 &  n_24090;
assign n_24093 = ~n_24091 & ~n_24092;
assign n_24094 =  x_2559 & ~n_24027;
assign n_24095 =  i_21 &  n_24027;
assign n_24096 = ~n_24094 & ~n_24095;
assign n_24097 =  x_2559 & ~n_24096;
assign n_24098 = ~x_2559 &  n_24096;
assign n_24099 = ~n_24097 & ~n_24098;
assign n_24100 =  x_2558 & ~n_24027;
assign n_24101 =  i_20 &  n_24027;
assign n_24102 = ~n_24100 & ~n_24101;
assign n_24103 =  x_2558 & ~n_24102;
assign n_24104 = ~x_2558 &  n_24102;
assign n_24105 = ~n_24103 & ~n_24104;
assign n_24106 =  x_2557 & ~n_24027;
assign n_24107 =  i_19 &  n_24027;
assign n_24108 = ~n_24106 & ~n_24107;
assign n_24109 =  x_2557 & ~n_24108;
assign n_24110 = ~x_2557 &  n_24108;
assign n_24111 = ~n_24109 & ~n_24110;
assign n_24112 =  x_2556 & ~n_24027;
assign n_24113 =  i_18 &  n_24027;
assign n_24114 = ~n_24112 & ~n_24113;
assign n_24115 =  x_2556 & ~n_24114;
assign n_24116 = ~x_2556 &  n_24114;
assign n_24117 = ~n_24115 & ~n_24116;
assign n_24118 =  x_2555 & ~n_24027;
assign n_24119 =  i_17 &  n_24027;
assign n_24120 = ~n_24118 & ~n_24119;
assign n_24121 =  x_2555 & ~n_24120;
assign n_24122 = ~x_2555 &  n_24120;
assign n_24123 = ~n_24121 & ~n_24122;
assign n_24124 =  x_2554 & ~n_24027;
assign n_24125 =  i_16 &  n_24027;
assign n_24126 = ~n_24124 & ~n_24125;
assign n_24127 =  x_2554 & ~n_24126;
assign n_24128 = ~x_2554 &  n_24126;
assign n_24129 = ~n_24127 & ~n_24128;
assign n_24130 =  x_2553 & ~n_24027;
assign n_24131 =  i_15 &  n_24027;
assign n_24132 = ~n_24130 & ~n_24131;
assign n_24133 =  x_2553 & ~n_24132;
assign n_24134 = ~x_2553 &  n_24132;
assign n_24135 = ~n_24133 & ~n_24134;
assign n_24136 =  x_2552 & ~n_24027;
assign n_24137 =  i_14 &  n_24027;
assign n_24138 = ~n_24136 & ~n_24137;
assign n_24139 =  x_2552 & ~n_24138;
assign n_24140 = ~x_2552 &  n_24138;
assign n_24141 = ~n_24139 & ~n_24140;
assign n_24142 =  x_2551 & ~n_24027;
assign n_24143 =  i_13 &  n_24027;
assign n_24144 = ~n_24142 & ~n_24143;
assign n_24145 =  x_2551 & ~n_24144;
assign n_24146 = ~x_2551 &  n_24144;
assign n_24147 = ~n_24145 & ~n_24146;
assign n_24148 =  x_2550 & ~n_24027;
assign n_24149 =  i_12 &  n_24027;
assign n_24150 = ~n_24148 & ~n_24149;
assign n_24151 =  x_2550 & ~n_24150;
assign n_24152 = ~x_2550 &  n_24150;
assign n_24153 = ~n_24151 & ~n_24152;
assign n_24154 =  x_2549 & ~n_24027;
assign n_24155 =  i_11 &  n_24027;
assign n_24156 = ~n_24154 & ~n_24155;
assign n_24157 =  x_2549 & ~n_24156;
assign n_24158 = ~x_2549 &  n_24156;
assign n_24159 = ~n_24157 & ~n_24158;
assign n_24160 =  x_2548 & ~n_24027;
assign n_24161 =  i_10 &  n_24027;
assign n_24162 = ~n_24160 & ~n_24161;
assign n_24163 =  x_2548 & ~n_24162;
assign n_24164 = ~x_2548 &  n_24162;
assign n_24165 = ~n_24163 & ~n_24164;
assign n_24166 =  x_2547 & ~n_24027;
assign n_24167 =  i_9 &  n_24027;
assign n_24168 = ~n_24166 & ~n_24167;
assign n_24169 =  x_2547 & ~n_24168;
assign n_24170 = ~x_2547 &  n_24168;
assign n_24171 = ~n_24169 & ~n_24170;
assign n_24172 =  x_2546 & ~n_24027;
assign n_24173 =  i_8 &  n_24027;
assign n_24174 = ~n_24172 & ~n_24173;
assign n_24175 =  x_2546 & ~n_24174;
assign n_24176 = ~x_2546 &  n_24174;
assign n_24177 = ~n_24175 & ~n_24176;
assign n_24178 =  x_2545 & ~n_24027;
assign n_24179 =  i_7 &  n_24027;
assign n_24180 = ~n_24178 & ~n_24179;
assign n_24181 =  x_2545 & ~n_24180;
assign n_24182 = ~x_2545 &  n_24180;
assign n_24183 = ~n_24181 & ~n_24182;
assign n_24184 =  x_2544 & ~n_24027;
assign n_24185 =  i_6 &  n_24027;
assign n_24186 = ~n_24184 & ~n_24185;
assign n_24187 =  x_2544 & ~n_24186;
assign n_24188 = ~x_2544 &  n_24186;
assign n_24189 = ~n_24187 & ~n_24188;
assign n_24190 =  x_2543 & ~n_24027;
assign n_24191 =  i_5 &  n_24027;
assign n_24192 = ~n_24190 & ~n_24191;
assign n_24193 =  x_2543 & ~n_24192;
assign n_24194 = ~x_2543 &  n_24192;
assign n_24195 = ~n_24193 & ~n_24194;
assign n_24196 =  x_2542 & ~n_24027;
assign n_24197 =  i_4 &  n_24027;
assign n_24198 = ~n_24196 & ~n_24197;
assign n_24199 =  x_2542 & ~n_24198;
assign n_24200 = ~x_2542 &  n_24198;
assign n_24201 = ~n_24199 & ~n_24200;
assign n_24202 =  x_2541 & ~n_24027;
assign n_24203 =  i_3 &  n_24027;
assign n_24204 = ~n_24202 & ~n_24203;
assign n_24205 =  x_2541 & ~n_24204;
assign n_24206 = ~x_2541 &  n_24204;
assign n_24207 = ~n_24205 & ~n_24206;
assign n_24208 =  x_2540 & ~n_24027;
assign n_24209 =  i_2 &  n_24027;
assign n_24210 = ~n_24208 & ~n_24209;
assign n_24211 =  x_2540 & ~n_24210;
assign n_24212 = ~x_2540 &  n_24210;
assign n_24213 = ~n_24211 & ~n_24212;
assign n_24214 =  x_2539 & ~n_24027;
assign n_24215 =  i_1 &  n_24027;
assign n_24216 = ~n_24214 & ~n_24215;
assign n_24217 =  x_2539 & ~n_24216;
assign n_24218 = ~x_2539 &  n_24216;
assign n_24219 = ~n_24217 & ~n_24218;
assign n_24220 =  n_1315 &  n_23892;
assign n_24221 =  x_2538 & ~n_24220;
assign n_24222 =  i_32 &  n_24220;
assign n_24223 = ~n_24221 & ~n_24222;
assign n_24224 =  x_2538 & ~n_24223;
assign n_24225 = ~x_2538 &  n_24223;
assign n_24226 = ~n_24224 & ~n_24225;
assign n_24227 =  x_2537 & ~n_24220;
assign n_24228 =  i_31 &  n_24220;
assign n_24229 = ~n_24227 & ~n_24228;
assign n_24230 =  x_2537 & ~n_24229;
assign n_24231 = ~x_2537 &  n_24229;
assign n_24232 = ~n_24230 & ~n_24231;
assign n_24233 =  x_2536 & ~n_24220;
assign n_24234 =  i_30 &  n_24220;
assign n_24235 = ~n_24233 & ~n_24234;
assign n_24236 =  x_2536 & ~n_24235;
assign n_24237 = ~x_2536 &  n_24235;
assign n_24238 = ~n_24236 & ~n_24237;
assign n_24239 =  x_2535 & ~n_24220;
assign n_24240 =  i_29 &  n_24220;
assign n_24241 = ~n_24239 & ~n_24240;
assign n_24242 =  x_2535 & ~n_24241;
assign n_24243 = ~x_2535 &  n_24241;
assign n_24244 = ~n_24242 & ~n_24243;
assign n_24245 =  x_2534 & ~n_24220;
assign n_24246 =  i_28 &  n_24220;
assign n_24247 = ~n_24245 & ~n_24246;
assign n_24248 =  x_2534 & ~n_24247;
assign n_24249 = ~x_2534 &  n_24247;
assign n_24250 = ~n_24248 & ~n_24249;
assign n_24251 =  x_2533 & ~n_24220;
assign n_24252 =  i_27 &  n_24220;
assign n_24253 = ~n_24251 & ~n_24252;
assign n_24254 =  x_2533 & ~n_24253;
assign n_24255 = ~x_2533 &  n_24253;
assign n_24256 = ~n_24254 & ~n_24255;
assign n_24257 =  x_2532 & ~n_24220;
assign n_24258 =  i_26 &  n_24220;
assign n_24259 = ~n_24257 & ~n_24258;
assign n_24260 =  x_2532 & ~n_24259;
assign n_24261 = ~x_2532 &  n_24259;
assign n_24262 = ~n_24260 & ~n_24261;
assign n_24263 =  x_2531 & ~n_24220;
assign n_24264 =  i_25 &  n_24220;
assign n_24265 = ~n_24263 & ~n_24264;
assign n_24266 =  x_2531 & ~n_24265;
assign n_24267 = ~x_2531 &  n_24265;
assign n_24268 = ~n_24266 & ~n_24267;
assign n_24269 =  x_2530 & ~n_24220;
assign n_24270 =  i_24 &  n_24220;
assign n_24271 = ~n_24269 & ~n_24270;
assign n_24272 =  x_2530 & ~n_24271;
assign n_24273 = ~x_2530 &  n_24271;
assign n_24274 = ~n_24272 & ~n_24273;
assign n_24275 =  x_2529 & ~n_24220;
assign n_24276 =  i_23 &  n_24220;
assign n_24277 = ~n_24275 & ~n_24276;
assign n_24278 =  x_2529 & ~n_24277;
assign n_24279 = ~x_2529 &  n_24277;
assign n_24280 = ~n_24278 & ~n_24279;
assign n_24281 =  x_2528 & ~n_24220;
assign n_24282 =  i_22 &  n_24220;
assign n_24283 = ~n_24281 & ~n_24282;
assign n_24284 =  x_2528 & ~n_24283;
assign n_24285 = ~x_2528 &  n_24283;
assign n_24286 = ~n_24284 & ~n_24285;
assign n_24287 =  x_2527 & ~n_24220;
assign n_24288 =  i_21 &  n_24220;
assign n_24289 = ~n_24287 & ~n_24288;
assign n_24290 =  x_2527 & ~n_24289;
assign n_24291 = ~x_2527 &  n_24289;
assign n_24292 = ~n_24290 & ~n_24291;
assign n_24293 =  x_2526 & ~n_24220;
assign n_24294 =  i_20 &  n_24220;
assign n_24295 = ~n_24293 & ~n_24294;
assign n_24296 =  x_2526 & ~n_24295;
assign n_24297 = ~x_2526 &  n_24295;
assign n_24298 = ~n_24296 & ~n_24297;
assign n_24299 =  x_2525 & ~n_24220;
assign n_24300 =  i_19 &  n_24220;
assign n_24301 = ~n_24299 & ~n_24300;
assign n_24302 =  x_2525 & ~n_24301;
assign n_24303 = ~x_2525 &  n_24301;
assign n_24304 = ~n_24302 & ~n_24303;
assign n_24305 =  x_2524 & ~n_24220;
assign n_24306 =  i_18 &  n_24220;
assign n_24307 = ~n_24305 & ~n_24306;
assign n_24308 =  x_2524 & ~n_24307;
assign n_24309 = ~x_2524 &  n_24307;
assign n_24310 = ~n_24308 & ~n_24309;
assign n_24311 =  x_2523 & ~n_24220;
assign n_24312 =  i_17 &  n_24220;
assign n_24313 = ~n_24311 & ~n_24312;
assign n_24314 =  x_2523 & ~n_24313;
assign n_24315 = ~x_2523 &  n_24313;
assign n_24316 = ~n_24314 & ~n_24315;
assign n_24317 =  x_2522 & ~n_24220;
assign n_24318 =  i_16 &  n_24220;
assign n_24319 = ~n_24317 & ~n_24318;
assign n_24320 =  x_2522 & ~n_24319;
assign n_24321 = ~x_2522 &  n_24319;
assign n_24322 = ~n_24320 & ~n_24321;
assign n_24323 =  x_2521 & ~n_24220;
assign n_24324 =  i_15 &  n_24220;
assign n_24325 = ~n_24323 & ~n_24324;
assign n_24326 =  x_2521 & ~n_24325;
assign n_24327 = ~x_2521 &  n_24325;
assign n_24328 = ~n_24326 & ~n_24327;
assign n_24329 =  x_2520 & ~n_24220;
assign n_24330 =  i_14 &  n_24220;
assign n_24331 = ~n_24329 & ~n_24330;
assign n_24332 =  x_2520 & ~n_24331;
assign n_24333 = ~x_2520 &  n_24331;
assign n_24334 = ~n_24332 & ~n_24333;
assign n_24335 =  x_2519 & ~n_24220;
assign n_24336 =  i_13 &  n_24220;
assign n_24337 = ~n_24335 & ~n_24336;
assign n_24338 =  x_2519 & ~n_24337;
assign n_24339 = ~x_2519 &  n_24337;
assign n_24340 = ~n_24338 & ~n_24339;
assign n_24341 =  x_2518 & ~n_24220;
assign n_24342 =  i_12 &  n_24220;
assign n_24343 = ~n_24341 & ~n_24342;
assign n_24344 =  x_2518 & ~n_24343;
assign n_24345 = ~x_2518 &  n_24343;
assign n_24346 = ~n_24344 & ~n_24345;
assign n_24347 =  x_2517 & ~n_24220;
assign n_24348 =  i_11 &  n_24220;
assign n_24349 = ~n_24347 & ~n_24348;
assign n_24350 =  x_2517 & ~n_24349;
assign n_24351 = ~x_2517 &  n_24349;
assign n_24352 = ~n_24350 & ~n_24351;
assign n_24353 =  x_2516 & ~n_24220;
assign n_24354 =  i_10 &  n_24220;
assign n_24355 = ~n_24353 & ~n_24354;
assign n_24356 =  x_2516 & ~n_24355;
assign n_24357 = ~x_2516 &  n_24355;
assign n_24358 = ~n_24356 & ~n_24357;
assign n_24359 =  x_2515 & ~n_24220;
assign n_24360 =  i_9 &  n_24220;
assign n_24361 = ~n_24359 & ~n_24360;
assign n_24362 =  x_2515 & ~n_24361;
assign n_24363 = ~x_2515 &  n_24361;
assign n_24364 = ~n_24362 & ~n_24363;
assign n_24365 =  x_2514 & ~n_24220;
assign n_24366 =  i_8 &  n_24220;
assign n_24367 = ~n_24365 & ~n_24366;
assign n_24368 =  x_2514 & ~n_24367;
assign n_24369 = ~x_2514 &  n_24367;
assign n_24370 = ~n_24368 & ~n_24369;
assign n_24371 =  x_2513 & ~n_24220;
assign n_24372 =  i_7 &  n_24220;
assign n_24373 = ~n_24371 & ~n_24372;
assign n_24374 =  x_2513 & ~n_24373;
assign n_24375 = ~x_2513 &  n_24373;
assign n_24376 = ~n_24374 & ~n_24375;
assign n_24377 =  x_2512 & ~n_24220;
assign n_24378 =  i_6 &  n_24220;
assign n_24379 = ~n_24377 & ~n_24378;
assign n_24380 =  x_2512 & ~n_24379;
assign n_24381 = ~x_2512 &  n_24379;
assign n_24382 = ~n_24380 & ~n_24381;
assign n_24383 =  x_2511 & ~n_24220;
assign n_24384 =  i_5 &  n_24220;
assign n_24385 = ~n_24383 & ~n_24384;
assign n_24386 =  x_2511 & ~n_24385;
assign n_24387 = ~x_2511 &  n_24385;
assign n_24388 = ~n_24386 & ~n_24387;
assign n_24389 =  x_2510 & ~n_24220;
assign n_24390 =  i_4 &  n_24220;
assign n_24391 = ~n_24389 & ~n_24390;
assign n_24392 =  x_2510 & ~n_24391;
assign n_24393 = ~x_2510 &  n_24391;
assign n_24394 = ~n_24392 & ~n_24393;
assign n_24395 =  x_2509 & ~n_24220;
assign n_24396 =  i_3 &  n_24220;
assign n_24397 = ~n_24395 & ~n_24396;
assign n_24398 =  x_2509 & ~n_24397;
assign n_24399 = ~x_2509 &  n_24397;
assign n_24400 = ~n_24398 & ~n_24399;
assign n_24401 =  x_2508 & ~n_24220;
assign n_24402 =  i_2 &  n_24220;
assign n_24403 = ~n_24401 & ~n_24402;
assign n_24404 =  x_2508 & ~n_24403;
assign n_24405 = ~x_2508 &  n_24403;
assign n_24406 = ~n_24404 & ~n_24405;
assign n_24407 =  x_2507 & ~n_24220;
assign n_24408 =  i_1 &  n_24220;
assign n_24409 = ~n_24407 & ~n_24408;
assign n_24410 =  x_2507 & ~n_24409;
assign n_24411 = ~x_2507 &  n_24409;
assign n_24412 = ~n_24410 & ~n_24411;
assign n_24413 =  n_389 &  n_980;
assign n_24414 =  n_982 &  n_24413;
assign n_24415 =  x_2506 & ~n_24414;
assign n_24416 =  i_32 &  n_24414;
assign n_24417 = ~n_24415 & ~n_24416;
assign n_24418 =  x_2506 & ~n_24417;
assign n_24419 = ~x_2506 &  n_24417;
assign n_24420 = ~n_24418 & ~n_24419;
assign n_24421 =  x_2505 & ~n_24414;
assign n_24422 =  i_31 &  n_24414;
assign n_24423 = ~n_24421 & ~n_24422;
assign n_24424 =  x_2505 & ~n_24423;
assign n_24425 = ~x_2505 &  n_24423;
assign n_24426 = ~n_24424 & ~n_24425;
assign n_24427 =  x_2504 & ~n_24414;
assign n_24428 =  i_30 &  n_24414;
assign n_24429 = ~n_24427 & ~n_24428;
assign n_24430 =  x_2504 & ~n_24429;
assign n_24431 = ~x_2504 &  n_24429;
assign n_24432 = ~n_24430 & ~n_24431;
assign n_24433 =  x_2503 & ~n_24414;
assign n_24434 =  i_29 &  n_24414;
assign n_24435 = ~n_24433 & ~n_24434;
assign n_24436 =  x_2503 & ~n_24435;
assign n_24437 = ~x_2503 &  n_24435;
assign n_24438 = ~n_24436 & ~n_24437;
assign n_24439 =  x_2502 & ~n_24414;
assign n_24440 =  i_28 &  n_24414;
assign n_24441 = ~n_24439 & ~n_24440;
assign n_24442 =  x_2502 & ~n_24441;
assign n_24443 = ~x_2502 &  n_24441;
assign n_24444 = ~n_24442 & ~n_24443;
assign n_24445 =  x_2501 & ~n_24414;
assign n_24446 =  i_27 &  n_24414;
assign n_24447 = ~n_24445 & ~n_24446;
assign n_24448 =  x_2501 & ~n_24447;
assign n_24449 = ~x_2501 &  n_24447;
assign n_24450 = ~n_24448 & ~n_24449;
assign n_24451 =  x_2500 & ~n_24414;
assign n_24452 =  i_26 &  n_24414;
assign n_24453 = ~n_24451 & ~n_24452;
assign n_24454 =  x_2500 & ~n_24453;
assign n_24455 = ~x_2500 &  n_24453;
assign n_24456 = ~n_24454 & ~n_24455;
assign n_24457 =  x_2499 & ~n_24414;
assign n_24458 =  i_25 &  n_24414;
assign n_24459 = ~n_24457 & ~n_24458;
assign n_24460 =  x_2499 & ~n_24459;
assign n_24461 = ~x_2499 &  n_24459;
assign n_24462 = ~n_24460 & ~n_24461;
assign n_24463 =  x_2498 & ~n_24414;
assign n_24464 =  i_24 &  n_24414;
assign n_24465 = ~n_24463 & ~n_24464;
assign n_24466 =  x_2498 & ~n_24465;
assign n_24467 = ~x_2498 &  n_24465;
assign n_24468 = ~n_24466 & ~n_24467;
assign n_24469 =  x_2497 & ~n_24414;
assign n_24470 =  i_23 &  n_24414;
assign n_24471 = ~n_24469 & ~n_24470;
assign n_24472 =  x_2497 & ~n_24471;
assign n_24473 = ~x_2497 &  n_24471;
assign n_24474 = ~n_24472 & ~n_24473;
assign n_24475 =  x_2496 & ~n_24414;
assign n_24476 =  i_22 &  n_24414;
assign n_24477 = ~n_24475 & ~n_24476;
assign n_24478 =  x_2496 & ~n_24477;
assign n_24479 = ~x_2496 &  n_24477;
assign n_24480 = ~n_24478 & ~n_24479;
assign n_24481 =  x_2495 & ~n_24414;
assign n_24482 =  i_21 &  n_24414;
assign n_24483 = ~n_24481 & ~n_24482;
assign n_24484 =  x_2495 & ~n_24483;
assign n_24485 = ~x_2495 &  n_24483;
assign n_24486 = ~n_24484 & ~n_24485;
assign n_24487 =  x_2494 & ~n_24414;
assign n_24488 =  i_20 &  n_24414;
assign n_24489 = ~n_24487 & ~n_24488;
assign n_24490 =  x_2494 & ~n_24489;
assign n_24491 = ~x_2494 &  n_24489;
assign n_24492 = ~n_24490 & ~n_24491;
assign n_24493 =  x_2493 & ~n_24414;
assign n_24494 =  i_19 &  n_24414;
assign n_24495 = ~n_24493 & ~n_24494;
assign n_24496 =  x_2493 & ~n_24495;
assign n_24497 = ~x_2493 &  n_24495;
assign n_24498 = ~n_24496 & ~n_24497;
assign n_24499 =  x_2492 & ~n_24414;
assign n_24500 =  i_18 &  n_24414;
assign n_24501 = ~n_24499 & ~n_24500;
assign n_24502 =  x_2492 & ~n_24501;
assign n_24503 = ~x_2492 &  n_24501;
assign n_24504 = ~n_24502 & ~n_24503;
assign n_24505 =  x_2491 & ~n_24414;
assign n_24506 =  i_17 &  n_24414;
assign n_24507 = ~n_24505 & ~n_24506;
assign n_24508 =  x_2491 & ~n_24507;
assign n_24509 = ~x_2491 &  n_24507;
assign n_24510 = ~n_24508 & ~n_24509;
assign n_24511 =  x_2490 & ~n_24414;
assign n_24512 =  i_16 &  n_24414;
assign n_24513 = ~n_24511 & ~n_24512;
assign n_24514 =  x_2490 & ~n_24513;
assign n_24515 = ~x_2490 &  n_24513;
assign n_24516 = ~n_24514 & ~n_24515;
assign n_24517 =  x_2489 & ~n_24414;
assign n_24518 =  i_15 &  n_24414;
assign n_24519 = ~n_24517 & ~n_24518;
assign n_24520 =  x_2489 & ~n_24519;
assign n_24521 = ~x_2489 &  n_24519;
assign n_24522 = ~n_24520 & ~n_24521;
assign n_24523 =  x_2488 & ~n_24414;
assign n_24524 =  i_14 &  n_24414;
assign n_24525 = ~n_24523 & ~n_24524;
assign n_24526 =  x_2488 & ~n_24525;
assign n_24527 = ~x_2488 &  n_24525;
assign n_24528 = ~n_24526 & ~n_24527;
assign n_24529 =  x_2487 & ~n_24414;
assign n_24530 =  i_13 &  n_24414;
assign n_24531 = ~n_24529 & ~n_24530;
assign n_24532 =  x_2487 & ~n_24531;
assign n_24533 = ~x_2487 &  n_24531;
assign n_24534 = ~n_24532 & ~n_24533;
assign n_24535 =  x_2486 & ~n_24414;
assign n_24536 =  i_12 &  n_24414;
assign n_24537 = ~n_24535 & ~n_24536;
assign n_24538 =  x_2486 & ~n_24537;
assign n_24539 = ~x_2486 &  n_24537;
assign n_24540 = ~n_24538 & ~n_24539;
assign n_24541 =  x_2485 & ~n_24414;
assign n_24542 =  i_11 &  n_24414;
assign n_24543 = ~n_24541 & ~n_24542;
assign n_24544 =  x_2485 & ~n_24543;
assign n_24545 = ~x_2485 &  n_24543;
assign n_24546 = ~n_24544 & ~n_24545;
assign n_24547 =  x_2484 & ~n_24414;
assign n_24548 =  i_10 &  n_24414;
assign n_24549 = ~n_24547 & ~n_24548;
assign n_24550 =  x_2484 & ~n_24549;
assign n_24551 = ~x_2484 &  n_24549;
assign n_24552 = ~n_24550 & ~n_24551;
assign n_24553 =  x_2483 & ~n_24414;
assign n_24554 =  i_9 &  n_24414;
assign n_24555 = ~n_24553 & ~n_24554;
assign n_24556 =  x_2483 & ~n_24555;
assign n_24557 = ~x_2483 &  n_24555;
assign n_24558 = ~n_24556 & ~n_24557;
assign n_24559 =  x_2482 & ~n_24414;
assign n_24560 =  i_8 &  n_24414;
assign n_24561 = ~n_24559 & ~n_24560;
assign n_24562 =  x_2482 & ~n_24561;
assign n_24563 = ~x_2482 &  n_24561;
assign n_24564 = ~n_24562 & ~n_24563;
assign n_24565 =  x_2481 & ~n_24414;
assign n_24566 =  i_7 &  n_24414;
assign n_24567 = ~n_24565 & ~n_24566;
assign n_24568 =  x_2481 & ~n_24567;
assign n_24569 = ~x_2481 &  n_24567;
assign n_24570 = ~n_24568 & ~n_24569;
assign n_24571 =  x_2480 & ~n_24414;
assign n_24572 =  i_6 &  n_24414;
assign n_24573 = ~n_24571 & ~n_24572;
assign n_24574 =  x_2480 & ~n_24573;
assign n_24575 = ~x_2480 &  n_24573;
assign n_24576 = ~n_24574 & ~n_24575;
assign n_24577 =  x_2479 & ~n_24414;
assign n_24578 =  i_5 &  n_24414;
assign n_24579 = ~n_24577 & ~n_24578;
assign n_24580 =  x_2479 & ~n_24579;
assign n_24581 = ~x_2479 &  n_24579;
assign n_24582 = ~n_24580 & ~n_24581;
assign n_24583 =  x_2478 & ~n_24414;
assign n_24584 =  i_4 &  n_24414;
assign n_24585 = ~n_24583 & ~n_24584;
assign n_24586 =  x_2478 & ~n_24585;
assign n_24587 = ~x_2478 &  n_24585;
assign n_24588 = ~n_24586 & ~n_24587;
assign n_24589 =  x_2477 & ~n_24414;
assign n_24590 =  i_3 &  n_24414;
assign n_24591 = ~n_24589 & ~n_24590;
assign n_24592 =  x_2477 & ~n_24591;
assign n_24593 = ~x_2477 &  n_24591;
assign n_24594 = ~n_24592 & ~n_24593;
assign n_24595 =  x_2476 & ~n_24414;
assign n_24596 =  i_2 &  n_24414;
assign n_24597 = ~n_24595 & ~n_24596;
assign n_24598 =  x_2476 & ~n_24597;
assign n_24599 = ~x_2476 &  n_24597;
assign n_24600 = ~n_24598 & ~n_24599;
assign n_24601 =  x_2475 & ~n_24414;
assign n_24602 =  i_1 &  n_24414;
assign n_24603 = ~n_24601 & ~n_24602;
assign n_24604 =  x_2475 & ~n_24603;
assign n_24605 = ~x_2475 &  n_24603;
assign n_24606 = ~n_24604 & ~n_24605;
assign n_24607 =  n_1 &  n_2303;
assign n_24608 = ~x_42 &  n_24607;
assign n_24609 =  x_2474 & ~n_24608;
assign n_24610 =  i_32 &  n_24608;
assign n_24611 = ~n_24609 & ~n_24610;
assign n_24612 =  x_2474 & ~n_24611;
assign n_24613 = ~x_2474 &  n_24611;
assign n_24614 = ~n_24612 & ~n_24613;
assign n_24615 =  x_2473 & ~n_24608;
assign n_24616 =  i_31 &  n_24608;
assign n_24617 = ~n_24615 & ~n_24616;
assign n_24618 =  x_2473 & ~n_24617;
assign n_24619 = ~x_2473 &  n_24617;
assign n_24620 = ~n_24618 & ~n_24619;
assign n_24621 =  x_2472 & ~n_24608;
assign n_24622 =  i_30 &  n_24608;
assign n_24623 = ~n_24621 & ~n_24622;
assign n_24624 =  x_2472 & ~n_24623;
assign n_24625 = ~x_2472 &  n_24623;
assign n_24626 = ~n_24624 & ~n_24625;
assign n_24627 =  x_2471 & ~n_24608;
assign n_24628 =  i_29 &  n_24608;
assign n_24629 = ~n_24627 & ~n_24628;
assign n_24630 =  x_2471 & ~n_24629;
assign n_24631 = ~x_2471 &  n_24629;
assign n_24632 = ~n_24630 & ~n_24631;
assign n_24633 =  x_2470 & ~n_24608;
assign n_24634 =  i_28 &  n_24608;
assign n_24635 = ~n_24633 & ~n_24634;
assign n_24636 =  x_2470 & ~n_24635;
assign n_24637 = ~x_2470 &  n_24635;
assign n_24638 = ~n_24636 & ~n_24637;
assign n_24639 =  x_2469 & ~n_24608;
assign n_24640 =  i_27 &  n_24608;
assign n_24641 = ~n_24639 & ~n_24640;
assign n_24642 =  x_2469 & ~n_24641;
assign n_24643 = ~x_2469 &  n_24641;
assign n_24644 = ~n_24642 & ~n_24643;
assign n_24645 =  x_2468 & ~n_24608;
assign n_24646 =  i_26 &  n_24608;
assign n_24647 = ~n_24645 & ~n_24646;
assign n_24648 =  x_2468 & ~n_24647;
assign n_24649 = ~x_2468 &  n_24647;
assign n_24650 = ~n_24648 & ~n_24649;
assign n_24651 =  x_2467 & ~n_24608;
assign n_24652 =  i_25 &  n_24608;
assign n_24653 = ~n_24651 & ~n_24652;
assign n_24654 =  x_2467 & ~n_24653;
assign n_24655 = ~x_2467 &  n_24653;
assign n_24656 = ~n_24654 & ~n_24655;
assign n_24657 =  x_2466 & ~n_24608;
assign n_24658 =  i_24 &  n_24608;
assign n_24659 = ~n_24657 & ~n_24658;
assign n_24660 =  x_2466 & ~n_24659;
assign n_24661 = ~x_2466 &  n_24659;
assign n_24662 = ~n_24660 & ~n_24661;
assign n_24663 =  x_2465 & ~n_24608;
assign n_24664 =  i_23 &  n_24608;
assign n_24665 = ~n_24663 & ~n_24664;
assign n_24666 =  x_2465 & ~n_24665;
assign n_24667 = ~x_2465 &  n_24665;
assign n_24668 = ~n_24666 & ~n_24667;
assign n_24669 =  x_2464 & ~n_24608;
assign n_24670 =  i_22 &  n_24608;
assign n_24671 = ~n_24669 & ~n_24670;
assign n_24672 =  x_2464 & ~n_24671;
assign n_24673 = ~x_2464 &  n_24671;
assign n_24674 = ~n_24672 & ~n_24673;
assign n_24675 =  x_2463 & ~n_24608;
assign n_24676 =  i_21 &  n_24608;
assign n_24677 = ~n_24675 & ~n_24676;
assign n_24678 =  x_2463 & ~n_24677;
assign n_24679 = ~x_2463 &  n_24677;
assign n_24680 = ~n_24678 & ~n_24679;
assign n_24681 =  x_2462 & ~n_24608;
assign n_24682 =  i_20 &  n_24608;
assign n_24683 = ~n_24681 & ~n_24682;
assign n_24684 =  x_2462 & ~n_24683;
assign n_24685 = ~x_2462 &  n_24683;
assign n_24686 = ~n_24684 & ~n_24685;
assign n_24687 =  x_2461 & ~n_24608;
assign n_24688 =  i_19 &  n_24608;
assign n_24689 = ~n_24687 & ~n_24688;
assign n_24690 =  x_2461 & ~n_24689;
assign n_24691 = ~x_2461 &  n_24689;
assign n_24692 = ~n_24690 & ~n_24691;
assign n_24693 =  x_2460 & ~n_24608;
assign n_24694 =  i_18 &  n_24608;
assign n_24695 = ~n_24693 & ~n_24694;
assign n_24696 =  x_2460 & ~n_24695;
assign n_24697 = ~x_2460 &  n_24695;
assign n_24698 = ~n_24696 & ~n_24697;
assign n_24699 =  x_2459 & ~n_24608;
assign n_24700 =  i_17 &  n_24608;
assign n_24701 = ~n_24699 & ~n_24700;
assign n_24702 =  x_2459 & ~n_24701;
assign n_24703 = ~x_2459 &  n_24701;
assign n_24704 = ~n_24702 & ~n_24703;
assign n_24705 =  x_2458 & ~n_24608;
assign n_24706 =  i_16 &  n_24608;
assign n_24707 = ~n_24705 & ~n_24706;
assign n_24708 =  x_2458 & ~n_24707;
assign n_24709 = ~x_2458 &  n_24707;
assign n_24710 = ~n_24708 & ~n_24709;
assign n_24711 =  x_2457 & ~n_24608;
assign n_24712 =  i_15 &  n_24608;
assign n_24713 = ~n_24711 & ~n_24712;
assign n_24714 =  x_2457 & ~n_24713;
assign n_24715 = ~x_2457 &  n_24713;
assign n_24716 = ~n_24714 & ~n_24715;
assign n_24717 =  x_2456 & ~n_24608;
assign n_24718 =  i_14 &  n_24608;
assign n_24719 = ~n_24717 & ~n_24718;
assign n_24720 =  x_2456 & ~n_24719;
assign n_24721 = ~x_2456 &  n_24719;
assign n_24722 = ~n_24720 & ~n_24721;
assign n_24723 =  x_2455 & ~n_24608;
assign n_24724 =  i_13 &  n_24608;
assign n_24725 = ~n_24723 & ~n_24724;
assign n_24726 =  x_2455 & ~n_24725;
assign n_24727 = ~x_2455 &  n_24725;
assign n_24728 = ~n_24726 & ~n_24727;
assign n_24729 =  x_2454 & ~n_24608;
assign n_24730 =  i_12 &  n_24608;
assign n_24731 = ~n_24729 & ~n_24730;
assign n_24732 =  x_2454 & ~n_24731;
assign n_24733 = ~x_2454 &  n_24731;
assign n_24734 = ~n_24732 & ~n_24733;
assign n_24735 =  x_2453 & ~n_24608;
assign n_24736 =  i_11 &  n_24608;
assign n_24737 = ~n_24735 & ~n_24736;
assign n_24738 =  x_2453 & ~n_24737;
assign n_24739 = ~x_2453 &  n_24737;
assign n_24740 = ~n_24738 & ~n_24739;
assign n_24741 =  x_2452 & ~n_24608;
assign n_24742 =  i_10 &  n_24608;
assign n_24743 = ~n_24741 & ~n_24742;
assign n_24744 =  x_2452 & ~n_24743;
assign n_24745 = ~x_2452 &  n_24743;
assign n_24746 = ~n_24744 & ~n_24745;
assign n_24747 =  x_2451 & ~n_24608;
assign n_24748 =  i_9 &  n_24608;
assign n_24749 = ~n_24747 & ~n_24748;
assign n_24750 =  x_2451 & ~n_24749;
assign n_24751 = ~x_2451 &  n_24749;
assign n_24752 = ~n_24750 & ~n_24751;
assign n_24753 =  x_2450 & ~n_24608;
assign n_24754 =  i_8 &  n_24608;
assign n_24755 = ~n_24753 & ~n_24754;
assign n_24756 =  x_2450 & ~n_24755;
assign n_24757 = ~x_2450 &  n_24755;
assign n_24758 = ~n_24756 & ~n_24757;
assign n_24759 =  x_2449 & ~n_24608;
assign n_24760 =  i_7 &  n_24608;
assign n_24761 = ~n_24759 & ~n_24760;
assign n_24762 =  x_2449 & ~n_24761;
assign n_24763 = ~x_2449 &  n_24761;
assign n_24764 = ~n_24762 & ~n_24763;
assign n_24765 =  x_2448 & ~n_24608;
assign n_24766 =  i_6 &  n_24608;
assign n_24767 = ~n_24765 & ~n_24766;
assign n_24768 =  x_2448 & ~n_24767;
assign n_24769 = ~x_2448 &  n_24767;
assign n_24770 = ~n_24768 & ~n_24769;
assign n_24771 =  x_2447 & ~n_24608;
assign n_24772 =  i_5 &  n_24608;
assign n_24773 = ~n_24771 & ~n_24772;
assign n_24774 =  x_2447 & ~n_24773;
assign n_24775 = ~x_2447 &  n_24773;
assign n_24776 = ~n_24774 & ~n_24775;
assign n_24777 =  x_2446 & ~n_24608;
assign n_24778 =  i_4 &  n_24608;
assign n_24779 = ~n_24777 & ~n_24778;
assign n_24780 =  x_2446 & ~n_24779;
assign n_24781 = ~x_2446 &  n_24779;
assign n_24782 = ~n_24780 & ~n_24781;
assign n_24783 =  x_2445 & ~n_24608;
assign n_24784 =  i_3 &  n_24608;
assign n_24785 = ~n_24783 & ~n_24784;
assign n_24786 =  x_2445 & ~n_24785;
assign n_24787 = ~x_2445 &  n_24785;
assign n_24788 = ~n_24786 & ~n_24787;
assign n_24789 =  x_2444 & ~n_24608;
assign n_24790 =  i_2 &  n_24608;
assign n_24791 = ~n_24789 & ~n_24790;
assign n_24792 =  x_2444 & ~n_24791;
assign n_24793 = ~x_2444 &  n_24791;
assign n_24794 = ~n_24792 & ~n_24793;
assign n_24795 =  x_2443 & ~n_24608;
assign n_24796 =  i_1 &  n_24608;
assign n_24797 = ~n_24795 & ~n_24796;
assign n_24798 =  x_2443 & ~n_24797;
assign n_24799 = ~x_2443 &  n_24797;
assign n_24800 = ~n_24798 & ~n_24799;
assign n_24801 =  n_2298 &  n_185;
assign n_24802 =  n_24801 &  n_983;
assign n_24803 =  x_2442 & ~n_24802;
assign n_24804 =  i_32 &  n_24802;
assign n_24805 = ~n_24803 & ~n_24804;
assign n_24806 =  x_2442 & ~n_24805;
assign n_24807 = ~x_2442 &  n_24805;
assign n_24808 = ~n_24806 & ~n_24807;
assign n_24809 =  x_2441 & ~n_24802;
assign n_24810 =  i_31 &  n_24802;
assign n_24811 = ~n_24809 & ~n_24810;
assign n_24812 =  x_2441 & ~n_24811;
assign n_24813 = ~x_2441 &  n_24811;
assign n_24814 = ~n_24812 & ~n_24813;
assign n_24815 =  x_2440 & ~n_24802;
assign n_24816 =  i_30 &  n_24802;
assign n_24817 = ~n_24815 & ~n_24816;
assign n_24818 =  x_2440 & ~n_24817;
assign n_24819 = ~x_2440 &  n_24817;
assign n_24820 = ~n_24818 & ~n_24819;
assign n_24821 =  x_2439 & ~n_24802;
assign n_24822 =  i_29 &  n_24802;
assign n_24823 = ~n_24821 & ~n_24822;
assign n_24824 =  x_2439 & ~n_24823;
assign n_24825 = ~x_2439 &  n_24823;
assign n_24826 = ~n_24824 & ~n_24825;
assign n_24827 =  x_2438 & ~n_24802;
assign n_24828 =  i_28 &  n_24802;
assign n_24829 = ~n_24827 & ~n_24828;
assign n_24830 =  x_2438 & ~n_24829;
assign n_24831 = ~x_2438 &  n_24829;
assign n_24832 = ~n_24830 & ~n_24831;
assign n_24833 =  x_2437 & ~n_24802;
assign n_24834 =  i_27 &  n_24802;
assign n_24835 = ~n_24833 & ~n_24834;
assign n_24836 =  x_2437 & ~n_24835;
assign n_24837 = ~x_2437 &  n_24835;
assign n_24838 = ~n_24836 & ~n_24837;
assign n_24839 =  x_2436 & ~n_24802;
assign n_24840 =  i_26 &  n_24802;
assign n_24841 = ~n_24839 & ~n_24840;
assign n_24842 =  x_2436 & ~n_24841;
assign n_24843 = ~x_2436 &  n_24841;
assign n_24844 = ~n_24842 & ~n_24843;
assign n_24845 =  x_2435 & ~n_24802;
assign n_24846 =  i_25 &  n_24802;
assign n_24847 = ~n_24845 & ~n_24846;
assign n_24848 =  x_2435 & ~n_24847;
assign n_24849 = ~x_2435 &  n_24847;
assign n_24850 = ~n_24848 & ~n_24849;
assign n_24851 =  x_2434 & ~n_24802;
assign n_24852 =  i_24 &  n_24802;
assign n_24853 = ~n_24851 & ~n_24852;
assign n_24854 =  x_2434 & ~n_24853;
assign n_24855 = ~x_2434 &  n_24853;
assign n_24856 = ~n_24854 & ~n_24855;
assign n_24857 =  x_2433 & ~n_24802;
assign n_24858 =  i_23 &  n_24802;
assign n_24859 = ~n_24857 & ~n_24858;
assign n_24860 =  x_2433 & ~n_24859;
assign n_24861 = ~x_2433 &  n_24859;
assign n_24862 = ~n_24860 & ~n_24861;
assign n_24863 =  x_2432 & ~n_24802;
assign n_24864 =  i_22 &  n_24802;
assign n_24865 = ~n_24863 & ~n_24864;
assign n_24866 =  x_2432 & ~n_24865;
assign n_24867 = ~x_2432 &  n_24865;
assign n_24868 = ~n_24866 & ~n_24867;
assign n_24869 =  x_2431 & ~n_24802;
assign n_24870 =  i_21 &  n_24802;
assign n_24871 = ~n_24869 & ~n_24870;
assign n_24872 =  x_2431 & ~n_24871;
assign n_24873 = ~x_2431 &  n_24871;
assign n_24874 = ~n_24872 & ~n_24873;
assign n_24875 =  x_2430 & ~n_24802;
assign n_24876 =  i_20 &  n_24802;
assign n_24877 = ~n_24875 & ~n_24876;
assign n_24878 =  x_2430 & ~n_24877;
assign n_24879 = ~x_2430 &  n_24877;
assign n_24880 = ~n_24878 & ~n_24879;
assign n_24881 =  x_2429 & ~n_24802;
assign n_24882 =  i_19 &  n_24802;
assign n_24883 = ~n_24881 & ~n_24882;
assign n_24884 =  x_2429 & ~n_24883;
assign n_24885 = ~x_2429 &  n_24883;
assign n_24886 = ~n_24884 & ~n_24885;
assign n_24887 =  x_2428 & ~n_24802;
assign n_24888 =  i_18 &  n_24802;
assign n_24889 = ~n_24887 & ~n_24888;
assign n_24890 =  x_2428 & ~n_24889;
assign n_24891 = ~x_2428 &  n_24889;
assign n_24892 = ~n_24890 & ~n_24891;
assign n_24893 =  x_2427 & ~n_24802;
assign n_24894 =  i_17 &  n_24802;
assign n_24895 = ~n_24893 & ~n_24894;
assign n_24896 =  x_2427 & ~n_24895;
assign n_24897 = ~x_2427 &  n_24895;
assign n_24898 = ~n_24896 & ~n_24897;
assign n_24899 =  x_2426 & ~n_24802;
assign n_24900 =  i_16 &  n_24802;
assign n_24901 = ~n_24899 & ~n_24900;
assign n_24902 =  x_2426 & ~n_24901;
assign n_24903 = ~x_2426 &  n_24901;
assign n_24904 = ~n_24902 & ~n_24903;
assign n_24905 =  x_2425 & ~n_24802;
assign n_24906 =  i_15 &  n_24802;
assign n_24907 = ~n_24905 & ~n_24906;
assign n_24908 =  x_2425 & ~n_24907;
assign n_24909 = ~x_2425 &  n_24907;
assign n_24910 = ~n_24908 & ~n_24909;
assign n_24911 =  x_2424 & ~n_24802;
assign n_24912 =  i_14 &  n_24802;
assign n_24913 = ~n_24911 & ~n_24912;
assign n_24914 =  x_2424 & ~n_24913;
assign n_24915 = ~x_2424 &  n_24913;
assign n_24916 = ~n_24914 & ~n_24915;
assign n_24917 =  x_2423 & ~n_24802;
assign n_24918 =  i_13 &  n_24802;
assign n_24919 = ~n_24917 & ~n_24918;
assign n_24920 =  x_2423 & ~n_24919;
assign n_24921 = ~x_2423 &  n_24919;
assign n_24922 = ~n_24920 & ~n_24921;
assign n_24923 =  x_2422 & ~n_24802;
assign n_24924 =  i_12 &  n_24802;
assign n_24925 = ~n_24923 & ~n_24924;
assign n_24926 =  x_2422 & ~n_24925;
assign n_24927 = ~x_2422 &  n_24925;
assign n_24928 = ~n_24926 & ~n_24927;
assign n_24929 =  x_2421 & ~n_24802;
assign n_24930 =  i_11 &  n_24802;
assign n_24931 = ~n_24929 & ~n_24930;
assign n_24932 =  x_2421 & ~n_24931;
assign n_24933 = ~x_2421 &  n_24931;
assign n_24934 = ~n_24932 & ~n_24933;
assign n_24935 =  x_2420 & ~n_24802;
assign n_24936 =  i_10 &  n_24802;
assign n_24937 = ~n_24935 & ~n_24936;
assign n_24938 =  x_2420 & ~n_24937;
assign n_24939 = ~x_2420 &  n_24937;
assign n_24940 = ~n_24938 & ~n_24939;
assign n_24941 =  x_2419 & ~n_24802;
assign n_24942 =  i_9 &  n_24802;
assign n_24943 = ~n_24941 & ~n_24942;
assign n_24944 =  x_2419 & ~n_24943;
assign n_24945 = ~x_2419 &  n_24943;
assign n_24946 = ~n_24944 & ~n_24945;
assign n_24947 =  x_2418 & ~n_24802;
assign n_24948 =  i_8 &  n_24802;
assign n_24949 = ~n_24947 & ~n_24948;
assign n_24950 =  x_2418 & ~n_24949;
assign n_24951 = ~x_2418 &  n_24949;
assign n_24952 = ~n_24950 & ~n_24951;
assign n_24953 =  x_2417 & ~n_24802;
assign n_24954 =  i_7 &  n_24802;
assign n_24955 = ~n_24953 & ~n_24954;
assign n_24956 =  x_2417 & ~n_24955;
assign n_24957 = ~x_2417 &  n_24955;
assign n_24958 = ~n_24956 & ~n_24957;
assign n_24959 =  x_2416 & ~n_24802;
assign n_24960 =  i_6 &  n_24802;
assign n_24961 = ~n_24959 & ~n_24960;
assign n_24962 =  x_2416 & ~n_24961;
assign n_24963 = ~x_2416 &  n_24961;
assign n_24964 = ~n_24962 & ~n_24963;
assign n_24965 =  x_2415 & ~n_24802;
assign n_24966 =  i_5 &  n_24802;
assign n_24967 = ~n_24965 & ~n_24966;
assign n_24968 =  x_2415 & ~n_24967;
assign n_24969 = ~x_2415 &  n_24967;
assign n_24970 = ~n_24968 & ~n_24969;
assign n_24971 =  x_2414 & ~n_24802;
assign n_24972 =  i_4 &  n_24802;
assign n_24973 = ~n_24971 & ~n_24972;
assign n_24974 =  x_2414 & ~n_24973;
assign n_24975 = ~x_2414 &  n_24973;
assign n_24976 = ~n_24974 & ~n_24975;
assign n_24977 =  x_2413 & ~n_24802;
assign n_24978 =  i_3 &  n_24802;
assign n_24979 = ~n_24977 & ~n_24978;
assign n_24980 =  x_2413 & ~n_24979;
assign n_24981 = ~x_2413 &  n_24979;
assign n_24982 = ~n_24980 & ~n_24981;
assign n_24983 =  x_2412 & ~n_24802;
assign n_24984 =  i_2 &  n_24802;
assign n_24985 = ~n_24983 & ~n_24984;
assign n_24986 =  x_2412 & ~n_24985;
assign n_24987 = ~x_2412 &  n_24985;
assign n_24988 = ~n_24986 & ~n_24987;
assign n_24989 =  x_2411 & ~n_24802;
assign n_24990 =  i_1 &  n_24802;
assign n_24991 = ~n_24989 & ~n_24990;
assign n_24992 =  x_2411 & ~n_24991;
assign n_24993 = ~x_2411 &  n_24991;
assign n_24994 = ~n_24992 & ~n_24993;
assign n_24995 =  n_784 &  n_2296;
assign n_24996 =  x_2410 & ~n_24995;
assign n_24997 =  i_32 &  n_24995;
assign n_24998 = ~n_24996 & ~n_24997;
assign n_24999 =  x_2410 & ~n_24998;
assign n_25000 = ~x_2410 &  n_24998;
assign n_25001 = ~n_24999 & ~n_25000;
assign n_25002 =  x_2409 & ~n_24995;
assign n_25003 =  i_31 &  n_24995;
assign n_25004 = ~n_25002 & ~n_25003;
assign n_25005 =  x_2409 & ~n_25004;
assign n_25006 = ~x_2409 &  n_25004;
assign n_25007 = ~n_25005 & ~n_25006;
assign n_25008 =  x_2408 & ~n_24995;
assign n_25009 =  i_30 &  n_24995;
assign n_25010 = ~n_25008 & ~n_25009;
assign n_25011 =  x_2408 & ~n_25010;
assign n_25012 = ~x_2408 &  n_25010;
assign n_25013 = ~n_25011 & ~n_25012;
assign n_25014 =  x_2407 & ~n_24995;
assign n_25015 =  i_29 &  n_24995;
assign n_25016 = ~n_25014 & ~n_25015;
assign n_25017 =  x_2407 & ~n_25016;
assign n_25018 = ~x_2407 &  n_25016;
assign n_25019 = ~n_25017 & ~n_25018;
assign n_25020 =  x_2406 & ~n_24995;
assign n_25021 =  i_28 &  n_24995;
assign n_25022 = ~n_25020 & ~n_25021;
assign n_25023 =  x_2406 & ~n_25022;
assign n_25024 = ~x_2406 &  n_25022;
assign n_25025 = ~n_25023 & ~n_25024;
assign n_25026 =  x_2405 & ~n_24995;
assign n_25027 =  i_27 &  n_24995;
assign n_25028 = ~n_25026 & ~n_25027;
assign n_25029 =  x_2405 & ~n_25028;
assign n_25030 = ~x_2405 &  n_25028;
assign n_25031 = ~n_25029 & ~n_25030;
assign n_25032 =  x_2404 & ~n_24995;
assign n_25033 =  i_26 &  n_24995;
assign n_25034 = ~n_25032 & ~n_25033;
assign n_25035 =  x_2404 & ~n_25034;
assign n_25036 = ~x_2404 &  n_25034;
assign n_25037 = ~n_25035 & ~n_25036;
assign n_25038 =  x_2403 & ~n_24995;
assign n_25039 =  i_25 &  n_24995;
assign n_25040 = ~n_25038 & ~n_25039;
assign n_25041 =  x_2403 & ~n_25040;
assign n_25042 = ~x_2403 &  n_25040;
assign n_25043 = ~n_25041 & ~n_25042;
assign n_25044 =  x_2402 & ~n_24995;
assign n_25045 =  i_24 &  n_24995;
assign n_25046 = ~n_25044 & ~n_25045;
assign n_25047 =  x_2402 & ~n_25046;
assign n_25048 = ~x_2402 &  n_25046;
assign n_25049 = ~n_25047 & ~n_25048;
assign n_25050 =  x_2401 & ~n_24995;
assign n_25051 =  i_23 &  n_24995;
assign n_25052 = ~n_25050 & ~n_25051;
assign n_25053 =  x_2401 & ~n_25052;
assign n_25054 = ~x_2401 &  n_25052;
assign n_25055 = ~n_25053 & ~n_25054;
assign n_25056 =  x_2400 & ~n_24995;
assign n_25057 =  i_22 &  n_24995;
assign n_25058 = ~n_25056 & ~n_25057;
assign n_25059 =  x_2400 & ~n_25058;
assign n_25060 = ~x_2400 &  n_25058;
assign n_25061 = ~n_25059 & ~n_25060;
assign n_25062 =  x_2399 & ~n_24995;
assign n_25063 =  i_21 &  n_24995;
assign n_25064 = ~n_25062 & ~n_25063;
assign n_25065 =  x_2399 & ~n_25064;
assign n_25066 = ~x_2399 &  n_25064;
assign n_25067 = ~n_25065 & ~n_25066;
assign n_25068 =  x_2398 & ~n_24995;
assign n_25069 =  i_20 &  n_24995;
assign n_25070 = ~n_25068 & ~n_25069;
assign n_25071 =  x_2398 & ~n_25070;
assign n_25072 = ~x_2398 &  n_25070;
assign n_25073 = ~n_25071 & ~n_25072;
assign n_25074 =  x_2397 & ~n_24995;
assign n_25075 =  i_19 &  n_24995;
assign n_25076 = ~n_25074 & ~n_25075;
assign n_25077 =  x_2397 & ~n_25076;
assign n_25078 = ~x_2397 &  n_25076;
assign n_25079 = ~n_25077 & ~n_25078;
assign n_25080 =  x_2396 & ~n_24995;
assign n_25081 =  i_18 &  n_24995;
assign n_25082 = ~n_25080 & ~n_25081;
assign n_25083 =  x_2396 & ~n_25082;
assign n_25084 = ~x_2396 &  n_25082;
assign n_25085 = ~n_25083 & ~n_25084;
assign n_25086 =  x_2395 & ~n_24995;
assign n_25087 =  i_17 &  n_24995;
assign n_25088 = ~n_25086 & ~n_25087;
assign n_25089 =  x_2395 & ~n_25088;
assign n_25090 = ~x_2395 &  n_25088;
assign n_25091 = ~n_25089 & ~n_25090;
assign n_25092 =  x_2394 & ~n_24995;
assign n_25093 =  i_16 &  n_24995;
assign n_25094 = ~n_25092 & ~n_25093;
assign n_25095 =  x_2394 & ~n_25094;
assign n_25096 = ~x_2394 &  n_25094;
assign n_25097 = ~n_25095 & ~n_25096;
assign n_25098 =  x_2393 & ~n_24995;
assign n_25099 =  i_15 &  n_24995;
assign n_25100 = ~n_25098 & ~n_25099;
assign n_25101 =  x_2393 & ~n_25100;
assign n_25102 = ~x_2393 &  n_25100;
assign n_25103 = ~n_25101 & ~n_25102;
assign n_25104 =  x_2392 & ~n_24995;
assign n_25105 =  i_14 &  n_24995;
assign n_25106 = ~n_25104 & ~n_25105;
assign n_25107 =  x_2392 & ~n_25106;
assign n_25108 = ~x_2392 &  n_25106;
assign n_25109 = ~n_25107 & ~n_25108;
assign n_25110 =  x_2391 & ~n_24995;
assign n_25111 =  i_13 &  n_24995;
assign n_25112 = ~n_25110 & ~n_25111;
assign n_25113 =  x_2391 & ~n_25112;
assign n_25114 = ~x_2391 &  n_25112;
assign n_25115 = ~n_25113 & ~n_25114;
assign n_25116 =  x_2390 & ~n_24995;
assign n_25117 =  i_12 &  n_24995;
assign n_25118 = ~n_25116 & ~n_25117;
assign n_25119 =  x_2390 & ~n_25118;
assign n_25120 = ~x_2390 &  n_25118;
assign n_25121 = ~n_25119 & ~n_25120;
assign n_25122 =  x_2389 & ~n_24995;
assign n_25123 =  i_11 &  n_24995;
assign n_25124 = ~n_25122 & ~n_25123;
assign n_25125 =  x_2389 & ~n_25124;
assign n_25126 = ~x_2389 &  n_25124;
assign n_25127 = ~n_25125 & ~n_25126;
assign n_25128 =  x_2388 & ~n_24995;
assign n_25129 =  i_10 &  n_24995;
assign n_25130 = ~n_25128 & ~n_25129;
assign n_25131 =  x_2388 & ~n_25130;
assign n_25132 = ~x_2388 &  n_25130;
assign n_25133 = ~n_25131 & ~n_25132;
assign n_25134 =  x_2387 & ~n_24995;
assign n_25135 =  i_9 &  n_24995;
assign n_25136 = ~n_25134 & ~n_25135;
assign n_25137 =  x_2387 & ~n_25136;
assign n_25138 = ~x_2387 &  n_25136;
assign n_25139 = ~n_25137 & ~n_25138;
assign n_25140 =  x_2386 & ~n_24995;
assign n_25141 =  i_8 &  n_24995;
assign n_25142 = ~n_25140 & ~n_25141;
assign n_25143 =  x_2386 & ~n_25142;
assign n_25144 = ~x_2386 &  n_25142;
assign n_25145 = ~n_25143 & ~n_25144;
assign n_25146 =  x_2385 & ~n_24995;
assign n_25147 =  i_7 &  n_24995;
assign n_25148 = ~n_25146 & ~n_25147;
assign n_25149 =  x_2385 & ~n_25148;
assign n_25150 = ~x_2385 &  n_25148;
assign n_25151 = ~n_25149 & ~n_25150;
assign n_25152 =  x_2384 & ~n_24995;
assign n_25153 =  i_6 &  n_24995;
assign n_25154 = ~n_25152 & ~n_25153;
assign n_25155 =  x_2384 & ~n_25154;
assign n_25156 = ~x_2384 &  n_25154;
assign n_25157 = ~n_25155 & ~n_25156;
assign n_25158 =  x_2383 & ~n_24995;
assign n_25159 =  i_5 &  n_24995;
assign n_25160 = ~n_25158 & ~n_25159;
assign n_25161 =  x_2383 & ~n_25160;
assign n_25162 = ~x_2383 &  n_25160;
assign n_25163 = ~n_25161 & ~n_25162;
assign n_25164 =  x_2382 & ~n_24995;
assign n_25165 =  i_4 &  n_24995;
assign n_25166 = ~n_25164 & ~n_25165;
assign n_25167 =  x_2382 & ~n_25166;
assign n_25168 = ~x_2382 &  n_25166;
assign n_25169 = ~n_25167 & ~n_25168;
assign n_25170 =  x_2381 & ~n_24995;
assign n_25171 =  i_3 &  n_24995;
assign n_25172 = ~n_25170 & ~n_25171;
assign n_25173 =  x_2381 & ~n_25172;
assign n_25174 = ~x_2381 &  n_25172;
assign n_25175 = ~n_25173 & ~n_25174;
assign n_25176 =  x_2380 & ~n_24995;
assign n_25177 =  i_2 &  n_24995;
assign n_25178 = ~n_25176 & ~n_25177;
assign n_25179 =  x_2380 & ~n_25178;
assign n_25180 = ~x_2380 &  n_25178;
assign n_25181 = ~n_25179 & ~n_25180;
assign n_25182 =  x_2379 & ~n_24995;
assign n_25183 =  i_1 &  n_24995;
assign n_25184 = ~n_25182 & ~n_25183;
assign n_25185 =  x_2379 & ~n_25184;
assign n_25186 = ~x_2379 &  n_25184;
assign n_25187 = ~n_25185 & ~n_25186;
assign n_25188 =  x_2378 & ~n_9;
assign n_25189 =  i_32 &  n_9;
assign n_25190 = ~n_25188 & ~n_25189;
assign n_25191 =  x_2378 & ~n_25190;
assign n_25192 = ~x_2378 &  n_25190;
assign n_25193 = ~n_25191 & ~n_25192;
assign n_25194 =  x_2377 & ~n_9;
assign n_25195 =  i_31 &  n_9;
assign n_25196 = ~n_25194 & ~n_25195;
assign n_25197 =  x_2377 & ~n_25196;
assign n_25198 = ~x_2377 &  n_25196;
assign n_25199 = ~n_25197 & ~n_25198;
assign n_25200 =  x_2376 & ~n_9;
assign n_25201 =  i_30 &  n_9;
assign n_25202 = ~n_25200 & ~n_25201;
assign n_25203 =  x_2376 & ~n_25202;
assign n_25204 = ~x_2376 &  n_25202;
assign n_25205 = ~n_25203 & ~n_25204;
assign n_25206 =  x_61 & ~n_22266;
assign n_25207 =  i_19 &  n_22266;
assign n_25208 = ~n_25206 & ~n_25207;
assign n_25209 =  x_61 & ~n_25208;
assign n_25210 = ~x_61 &  n_25208;
assign n_25211 = ~n_25209 & ~n_25210;
assign n_25212 =  x_60 & ~n_22266;
assign n_25213 =  i_18 &  n_22266;
assign n_25214 = ~n_25212 & ~n_25213;
assign n_25215 =  x_60 & ~n_25214;
assign n_25216 = ~x_60 &  n_25214;
assign n_25217 = ~n_25215 & ~n_25216;
assign n_25218 =  x_59 & ~n_22266;
assign n_25219 =  i_17 &  n_22266;
assign n_25220 = ~n_25218 & ~n_25219;
assign n_25221 =  x_59 & ~n_25220;
assign n_25222 = ~x_59 &  n_25220;
assign n_25223 = ~n_25221 & ~n_25222;
assign n_25224 =  x_58 & ~n_22266;
assign n_25225 =  i_16 &  n_22266;
assign n_25226 = ~n_25224 & ~n_25225;
assign n_25227 =  x_58 & ~n_25226;
assign n_25228 = ~x_58 &  n_25226;
assign n_25229 = ~n_25227 & ~n_25228;
assign n_25230 =  x_57 & ~n_22266;
assign n_25231 =  i_15 &  n_22266;
assign n_25232 = ~n_25230 & ~n_25231;
assign n_25233 =  x_57 & ~n_25232;
assign n_25234 = ~x_57 &  n_25232;
assign n_25235 = ~n_25233 & ~n_25234;
assign n_25236 =  x_56 & ~n_22266;
assign n_25237 =  i_14 &  n_22266;
assign n_25238 = ~n_25236 & ~n_25237;
assign n_25239 =  x_56 & ~n_25238;
assign n_25240 = ~x_56 &  n_25238;
assign n_25241 = ~n_25239 & ~n_25240;
assign n_25242 =  x_55 & ~n_22266;
assign n_25243 =  i_13 &  n_22266;
assign n_25244 = ~n_25242 & ~n_25243;
assign n_25245 =  x_55 & ~n_25244;
assign n_25246 = ~x_55 &  n_25244;
assign n_25247 = ~n_25245 & ~n_25246;
assign n_25248 =  x_54 & ~n_22266;
assign n_25249 =  i_12 &  n_22266;
assign n_25250 = ~n_25248 & ~n_25249;
assign n_25251 =  x_54 & ~n_25250;
assign n_25252 = ~x_54 &  n_25250;
assign n_25253 = ~n_25251 & ~n_25252;
assign n_25254 =  x_53 & ~n_22266;
assign n_25255 =  i_11 &  n_22266;
assign n_25256 = ~n_25254 & ~n_25255;
assign n_25257 =  x_53 & ~n_25256;
assign n_25258 = ~x_53 &  n_25256;
assign n_25259 = ~n_25257 & ~n_25258;
assign n_25260 =  x_52 & ~n_22266;
assign n_25261 =  i_10 &  n_22266;
assign n_25262 = ~n_25260 & ~n_25261;
assign n_25263 =  x_52 & ~n_25262;
assign n_25264 = ~x_52 &  n_25262;
assign n_25265 = ~n_25263 & ~n_25264;
assign n_25266 =  x_51 & ~n_22266;
assign n_25267 =  i_9 &  n_22266;
assign n_25268 = ~n_25266 & ~n_25267;
assign n_25269 =  x_51 & ~n_25268;
assign n_25270 = ~x_51 &  n_25268;
assign n_25271 = ~n_25269 & ~n_25270;
assign n_25272 =  x_50 & ~n_22266;
assign n_25273 =  i_8 &  n_22266;
assign n_25274 = ~n_25272 & ~n_25273;
assign n_25275 =  x_50 & ~n_25274;
assign n_25276 = ~x_50 &  n_25274;
assign n_25277 = ~n_25275 & ~n_25276;
assign n_25278 =  x_49 & ~n_22266;
assign n_25279 =  i_7 &  n_22266;
assign n_25280 = ~n_25278 & ~n_25279;
assign n_25281 =  x_49 & ~n_25280;
assign n_25282 = ~x_49 &  n_25280;
assign n_25283 = ~n_25281 & ~n_25282;
assign n_25284 =  x_48 & ~n_22266;
assign n_25285 =  i_6 &  n_22266;
assign n_25286 = ~n_25284 & ~n_25285;
assign n_25287 =  x_48 & ~n_25286;
assign n_25288 = ~x_48 &  n_25286;
assign n_25289 = ~n_25287 & ~n_25288;
assign n_25290 =  x_47 & ~n_22266;
assign n_25291 =  i_5 &  n_22266;
assign n_25292 = ~n_25290 & ~n_25291;
assign n_25293 =  x_47 & ~n_25292;
assign n_25294 = ~x_47 &  n_25292;
assign n_25295 = ~n_25293 & ~n_25294;
assign n_25296 =  x_46 & ~n_22266;
assign n_25297 =  i_4 &  n_22266;
assign n_25298 = ~n_25296 & ~n_25297;
assign n_25299 =  x_46 & ~n_25298;
assign n_25300 = ~x_46 &  n_25298;
assign n_25301 = ~n_25299 & ~n_25300;
assign n_25302 =  x_45 & ~n_22266;
assign n_25303 =  i_3 &  n_22266;
assign n_25304 = ~n_25302 & ~n_25303;
assign n_25305 =  x_45 & ~n_25304;
assign n_25306 = ~x_45 &  n_25304;
assign n_25307 = ~n_25305 & ~n_25306;
assign n_25308 =  x_44 & ~n_22266;
assign n_25309 =  i_2 &  n_22266;
assign n_25310 = ~n_25308 & ~n_25309;
assign n_25311 =  x_44 & ~n_25310;
assign n_25312 = ~x_44 &  n_25310;
assign n_25313 = ~n_25311 & ~n_25312;
assign n_25314 =  x_43 & ~n_22266;
assign n_25315 =  i_1 &  n_22266;
assign n_25316 = ~n_25314 & ~n_25315;
assign n_25317 =  x_43 & ~n_25316;
assign n_25318 = ~x_43 &  n_25316;
assign n_25319 = ~n_25317 & ~n_25318;
assign n_25320 =  n_1906 &  n_1179;
assign n_25321 = ~x_1608 & ~x_1609;
assign n_25322 = ~x_1607 &  n_25321;
assign n_25323 = ~x_1606 &  n_25322;
assign n_25324 = ~x_1605 & ~x_1610;
assign n_25325 =  n_25323 &  n_25324;
assign n_25326 = ~x_1604 &  n_25325;
assign n_25327 = ~x_1603 &  n_25326;
assign n_25328 = ~x_1602 &  n_25327;
assign n_25329 = ~x_1601 &  n_25328;
assign n_25330 = ~x_1600 &  n_25329;
assign n_25331 = ~x_1599 &  n_25330;
assign n_25332 = ~x_1598 &  n_25331;
assign n_25333 = ~x_1597 &  n_25332;
assign n_25334 = ~x_1596 &  n_25333;
assign n_25335 = ~x_1595 &  n_25334;
assign n_25336 = ~x_1594 &  n_25335;
assign n_25337 = ~x_1593 &  n_25336;
assign n_25338 = ~x_1592 &  n_25337;
assign n_25339 = ~x_1591 &  n_25338;
assign n_25340 = ~x_1590 &  n_25339;
assign n_25341 = ~x_1589 &  n_25340;
assign n_25342 = ~x_1588 &  n_25341;
assign n_25343 = ~x_1587 &  n_25342;
assign n_25344 = ~x_1586 &  n_25343;
assign n_25345 = ~x_1585 &  n_25344;
assign n_25346 = ~x_1584 &  n_25345;
assign n_25347 = ~x_1583 &  n_25346;
assign n_25348 = ~x_1582 &  n_25347;
assign n_25349 = ~x_1581 &  n_25348;
assign n_25350 =  x_1581 & ~n_25348;
assign n_25351 = ~n_25349 & ~n_25350;
assign n_25352 =  x_1583 & ~n_25346;
assign n_25353 = ~n_25347 & ~n_25352;
assign n_25354 =  x_1585 & ~n_25344;
assign n_25355 = ~n_25345 & ~n_25354;
assign n_25356 =  x_1587 & ~n_25342;
assign n_25357 = ~n_25343 & ~n_25356;
assign n_25358 =  x_1589 & ~n_25340;
assign n_25359 = ~n_25341 & ~n_25358;
assign n_25360 =  x_1591 & ~n_25338;
assign n_25361 = ~n_25339 & ~n_25360;
assign n_25362 =  x_1593 & ~n_25336;
assign n_25363 = ~n_25337 & ~n_25362;
assign n_25364 =  x_1595 & ~n_25334;
assign n_25365 = ~n_25335 & ~n_25364;
assign n_25366 =  x_1597 & ~n_25332;
assign n_25367 = ~n_25333 & ~n_25366;
assign n_25368 =  x_1599 & ~n_25330;
assign n_25369 = ~n_25331 & ~n_25368;
assign n_25370 =  x_1601 & ~n_25328;
assign n_25371 = ~n_25329 & ~n_25370;
assign n_25372 =  x_1603 & ~n_25326;
assign n_25373 = ~n_25327 & ~n_25372;
assign n_25374 = ~x_1605 &  x_1610;
assign n_25375 =  n_25323 &  n_25374;
assign n_25376 = ~x_1604 &  n_25375;
assign n_25377 =  n_25373 &  n_25376;
assign n_25378 = ~x_1602 &  n_25377;
assign n_25379 =  n_25371 &  n_25378;
assign n_25380 = ~x_1600 &  n_25379;
assign n_25381 =  n_25369 &  n_25380;
assign n_25382 = ~x_1598 &  n_25381;
assign n_25383 =  n_25367 &  n_25382;
assign n_25384 = ~x_1596 &  n_25383;
assign n_25385 =  n_25365 &  n_25384;
assign n_25386 = ~x_1594 &  n_25385;
assign n_25387 =  n_25363 &  n_25386;
assign n_25388 = ~x_1592 &  n_25387;
assign n_25389 =  n_25361 &  n_25388;
assign n_25390 = ~x_1590 &  n_25389;
assign n_25391 =  n_25359 &  n_25390;
assign n_25392 = ~x_1588 &  n_25391;
assign n_25393 =  n_25357 &  n_25392;
assign n_25394 = ~x_1586 &  n_25393;
assign n_25395 =  n_25355 &  n_25394;
assign n_25396 = ~x_1584 &  n_25395;
assign n_25397 =  n_25353 &  n_25396;
assign n_25398 = ~x_1582 &  n_25397;
assign n_25399 =  n_25351 &  n_25398;
assign n_25400 = ~x_1580 &  n_25399;
assign n_25401 = ~x_1580 &  n_25349;
assign n_25402 =  x_1580 & ~n_25349;
assign n_25403 = ~n_25401 & ~n_25402;
assign n_25404 = ~n_25399 & ~n_25403;
assign n_25405 = ~n_25400 & ~n_25404;
assign n_25406 = ~n_25351 & ~n_25398;
assign n_25407 = ~n_25399 & ~n_25406;
assign n_25408 =  x_1582 & ~n_25347;
assign n_25409 = ~n_25348 & ~n_25408;
assign n_25410 = ~n_25397 & ~n_25409;
assign n_25411 = ~n_25398 & ~n_25410;
assign n_25412 = ~n_25353 & ~n_25396;
assign n_25413 = ~n_25397 & ~n_25412;
assign n_25414 =  x_1584 & ~n_25345;
assign n_25415 = ~n_25346 & ~n_25414;
assign n_25416 = ~n_25395 & ~n_25415;
assign n_25417 = ~n_25396 & ~n_25416;
assign n_25418 = ~n_25355 & ~n_25394;
assign n_25419 = ~n_25395 & ~n_25418;
assign n_25420 =  x_1586 & ~n_25343;
assign n_25421 = ~n_25344 & ~n_25420;
assign n_25422 = ~n_25393 & ~n_25421;
assign n_25423 = ~n_25394 & ~n_25422;
assign n_25424 = ~n_25357 & ~n_25392;
assign n_25425 = ~n_25393 & ~n_25424;
assign n_25426 =  x_1588 & ~n_25341;
assign n_25427 = ~n_25342 & ~n_25426;
assign n_25428 = ~n_25391 & ~n_25427;
assign n_25429 = ~n_25392 & ~n_25428;
assign n_25430 = ~n_25359 & ~n_25390;
assign n_25431 = ~n_25391 & ~n_25430;
assign n_25432 =  x_1590 & ~n_25339;
assign n_25433 = ~n_25340 & ~n_25432;
assign n_25434 = ~n_25389 & ~n_25433;
assign n_25435 = ~n_25390 & ~n_25434;
assign n_25436 = ~n_25361 & ~n_25388;
assign n_25437 = ~n_25389 & ~n_25436;
assign n_25438 =  x_1592 & ~n_25337;
assign n_25439 = ~n_25338 & ~n_25438;
assign n_25440 = ~n_25387 & ~n_25439;
assign n_25441 = ~n_25388 & ~n_25440;
assign n_25442 = ~n_25363 & ~n_25386;
assign n_25443 = ~n_25387 & ~n_25442;
assign n_25444 =  x_1594 & ~n_25335;
assign n_25445 = ~n_25336 & ~n_25444;
assign n_25446 = ~n_25385 & ~n_25445;
assign n_25447 = ~n_25386 & ~n_25446;
assign n_25448 = ~n_25365 & ~n_25384;
assign n_25449 = ~n_25385 & ~n_25448;
assign n_25450 =  x_1596 & ~n_25333;
assign n_25451 = ~n_25334 & ~n_25450;
assign n_25452 = ~n_25383 & ~n_25451;
assign n_25453 = ~n_25384 & ~n_25452;
assign n_25454 = ~n_25367 & ~n_25382;
assign n_25455 = ~n_25383 & ~n_25454;
assign n_25456 =  x_1598 & ~n_25331;
assign n_25457 = ~n_25332 & ~n_25456;
assign n_25458 = ~n_25381 & ~n_25457;
assign n_25459 = ~n_25382 & ~n_25458;
assign n_25460 = ~n_25369 & ~n_25380;
assign n_25461 = ~n_25381 & ~n_25460;
assign n_25462 =  x_1600 & ~n_25329;
assign n_25463 = ~n_25330 & ~n_25462;
assign n_25464 = ~n_25379 & ~n_25463;
assign n_25465 = ~n_25380 & ~n_25464;
assign n_25466 = ~n_25371 & ~n_25378;
assign n_25467 = ~n_25379 & ~n_25466;
assign n_25468 =  x_1602 & ~n_25327;
assign n_25469 = ~n_25328 & ~n_25468;
assign n_25470 = ~n_25377 & ~n_25469;
assign n_25471 = ~n_25378 & ~n_25470;
assign n_25472 = ~n_25373 & ~n_25376;
assign n_25473 = ~n_25377 & ~n_25472;
assign n_25474 = ~n_25325 & ~n_25375;
assign n_25475 =  x_1604 & ~n_25474;
assign n_25476 = ~x_1604 &  n_25474;
assign n_25477 = ~n_25475 & ~n_25476;
assign n_25478 =  x_1605 & ~n_25323;
assign n_25479 =  n_25474 & ~n_25478;
assign n_25480 =  x_1607 & ~n_25321;
assign n_25481 = ~n_25322 & ~n_25480;
assign n_25482 = ~x_1545 & ~x_1609;
assign n_25483 =  x_1546 & ~x_1610;
assign n_25484 =  x_1545 &  x_1609;
assign n_25485 = ~n_25483 & ~n_25484;
assign n_25486 = ~n_25482 & ~n_25485;
assign n_25487 = ~x_1544 & ~n_25486;
assign n_25488 =  x_1544 &  n_25486;
assign n_25489 =  x_1608 & ~x_1609;
assign n_25490 = ~x_1608 &  x_1609;
assign n_25491 = ~n_25489 & ~n_25490;
assign n_25492 = ~n_25488 &  n_25491;
assign n_25493 = ~n_25487 & ~n_25492;
assign n_25494 = ~n_25481 & ~n_25493;
assign n_25495 =  n_25481 &  n_25493;
assign n_25496 = ~x_1543 & ~n_25495;
assign n_25497 = ~n_25494 & ~n_25496;
assign n_25498 =  x_1606 & ~n_25322;
assign n_25499 = ~n_25323 & ~n_25498;
assign n_25500 = ~n_25497 & ~n_25499;
assign n_25501 =  n_25497 &  n_25499;
assign n_25502 = ~x_1542 & ~n_25501;
assign n_25503 = ~n_25500 & ~n_25502;
assign n_25504 = ~n_25479 & ~n_25503;
assign n_25505 =  n_25479 &  n_25503;
assign n_25506 = ~x_1541 & ~n_25505;
assign n_25507 = ~n_25504 & ~n_25506;
assign n_25508 =  n_25477 & ~n_25507;
assign n_25509 = ~n_25477 &  n_25507;
assign n_25510 = ~x_1540 & ~n_25509;
assign n_25511 = ~n_25508 & ~n_25510;
assign n_25512 = ~n_25473 & ~n_25511;
assign n_25513 =  n_25473 &  n_25511;
assign n_25514 = ~x_1539 & ~n_25513;
assign n_25515 = ~n_25512 & ~n_25514;
assign n_25516 = ~n_25471 & ~n_25515;
assign n_25517 =  n_25471 &  n_25515;
assign n_25518 = ~x_1538 & ~n_25517;
assign n_25519 = ~n_25516 & ~n_25518;
assign n_25520 = ~n_25467 & ~n_25519;
assign n_25521 =  n_25467 &  n_25519;
assign n_25522 = ~x_1537 & ~n_25521;
assign n_25523 = ~n_25520 & ~n_25522;
assign n_25524 = ~n_25465 & ~n_25523;
assign n_25525 =  n_25465 &  n_25523;
assign n_25526 = ~x_1536 & ~n_25525;
assign n_25527 = ~n_25524 & ~n_25526;
assign n_25528 = ~n_25461 & ~n_25527;
assign n_25529 =  n_25461 &  n_25527;
assign n_25530 = ~x_1535 & ~n_25529;
assign n_25531 = ~n_25528 & ~n_25530;
assign n_25532 = ~n_25459 & ~n_25531;
assign n_25533 =  n_25459 &  n_25531;
assign n_25534 = ~x_1534 & ~n_25533;
assign n_25535 = ~n_25532 & ~n_25534;
assign n_25536 = ~n_25455 & ~n_25535;
assign n_25537 =  n_25455 &  n_25535;
assign n_25538 = ~x_1533 & ~n_25537;
assign n_25539 = ~n_25536 & ~n_25538;
assign n_25540 = ~n_25453 & ~n_25539;
assign n_25541 =  n_25453 &  n_25539;
assign n_25542 = ~x_1532 & ~n_25541;
assign n_25543 = ~n_25540 & ~n_25542;
assign n_25544 = ~n_25449 & ~n_25543;
assign n_25545 =  n_25449 &  n_25543;
assign n_25546 = ~x_1531 & ~n_25545;
assign n_25547 = ~n_25544 & ~n_25546;
assign n_25548 = ~n_25447 & ~n_25547;
assign n_25549 =  n_25447 &  n_25547;
assign n_25550 = ~x_1530 & ~n_25549;
assign n_25551 = ~n_25548 & ~n_25550;
assign n_25552 = ~n_25443 & ~n_25551;
assign n_25553 =  n_25443 &  n_25551;
assign n_25554 = ~x_1529 & ~n_25553;
assign n_25555 = ~n_25552 & ~n_25554;
assign n_25556 = ~n_25441 & ~n_25555;
assign n_25557 =  n_25441 &  n_25555;
assign n_25558 = ~x_1528 & ~n_25557;
assign n_25559 = ~n_25556 & ~n_25558;
assign n_25560 = ~n_25437 & ~n_25559;
assign n_25561 =  n_25437 &  n_25559;
assign n_25562 = ~x_1527 & ~n_25561;
assign n_25563 = ~n_25560 & ~n_25562;
assign n_25564 = ~n_25435 & ~n_25563;
assign n_25565 =  n_25435 &  n_25563;
assign n_25566 = ~x_1526 & ~n_25565;
assign n_25567 = ~n_25564 & ~n_25566;
assign n_25568 = ~n_25431 & ~n_25567;
assign n_25569 =  n_25431 &  n_25567;
assign n_25570 = ~x_1525 & ~n_25569;
assign n_25571 = ~n_25568 & ~n_25570;
assign n_25572 = ~n_25429 & ~n_25571;
assign n_25573 =  n_25429 &  n_25571;
assign n_25574 = ~x_1524 & ~n_25573;
assign n_25575 = ~n_25572 & ~n_25574;
assign n_25576 = ~n_25425 & ~n_25575;
assign n_25577 =  n_25425 &  n_25575;
assign n_25578 = ~x_1523 & ~n_25577;
assign n_25579 = ~n_25576 & ~n_25578;
assign n_25580 = ~n_25423 & ~n_25579;
assign n_25581 =  n_25423 &  n_25579;
assign n_25582 = ~x_1522 & ~n_25581;
assign n_25583 = ~n_25580 & ~n_25582;
assign n_25584 = ~n_25419 & ~n_25583;
assign n_25585 =  n_25419 &  n_25583;
assign n_25586 = ~x_1521 & ~n_25585;
assign n_25587 = ~n_25584 & ~n_25586;
assign n_25588 = ~n_25417 & ~n_25587;
assign n_25589 =  n_25417 &  n_25587;
assign n_25590 = ~x_1520 & ~n_25589;
assign n_25591 = ~n_25588 & ~n_25590;
assign n_25592 = ~n_25413 & ~n_25591;
assign n_25593 =  n_25413 &  n_25591;
assign n_25594 = ~x_1519 & ~n_25593;
assign n_25595 = ~n_25592 & ~n_25594;
assign n_25596 = ~n_25411 & ~n_25595;
assign n_25597 =  n_25411 &  n_25595;
assign n_25598 = ~x_1518 & ~n_25597;
assign n_25599 = ~n_25596 & ~n_25598;
assign n_25600 = ~n_25407 & ~n_25599;
assign n_25601 =  n_25407 &  n_25599;
assign n_25602 = ~x_1517 & ~n_25601;
assign n_25603 = ~n_25600 & ~n_25602;
assign n_25604 = ~n_25405 & ~n_25603;
assign n_25605 =  n_25405 &  n_25603;
assign n_25606 = ~n_25604 & ~n_25605;
assign n_25607 = ~x_1516 & ~n_25606;
assign n_25608 =  x_1516 &  n_25606;
assign n_25609 = ~n_25607 & ~n_25608;
assign n_25610 = ~x_1579 & ~n_25401;
assign n_25611 = ~n_25400 &  n_25610;
assign n_25612 = ~x_1516 & ~n_25605;
assign n_25613 = ~n_25604 & ~n_25612;
assign n_25614 =  n_25611 & ~n_25613;
assign n_25615 = ~n_25600 & ~n_25601;
assign n_25616 =  x_1517 &  n_25615;
assign n_25617 = ~x_1517 & ~n_25615;
assign n_25618 = ~n_25616 & ~n_25617;
assign n_25619 = ~n_25596 & ~n_25597;
assign n_25620 =  x_1518 &  n_25619;
assign n_25621 = ~x_1518 & ~n_25619;
assign n_25622 = ~n_25620 & ~n_25621;
assign n_25623 = ~n_25592 & ~n_25593;
assign n_25624 =  x_1519 &  n_25623;
assign n_25625 = ~x_1519 & ~n_25623;
assign n_25626 = ~n_25624 & ~n_25625;
assign n_25627 = ~n_25588 & ~n_25589;
assign n_25628 =  x_1520 &  n_25627;
assign n_25629 = ~x_1520 & ~n_25627;
assign n_25630 = ~n_25628 & ~n_25629;
assign n_25631 = ~n_25584 & ~n_25585;
assign n_25632 =  x_1521 &  n_25631;
assign n_25633 = ~x_1521 & ~n_25631;
assign n_25634 = ~n_25632 & ~n_25633;
assign n_25635 = ~n_25580 & ~n_25581;
assign n_25636 =  x_1522 &  n_25635;
assign n_25637 = ~x_1522 & ~n_25635;
assign n_25638 = ~n_25636 & ~n_25637;
assign n_25639 = ~n_25576 & ~n_25577;
assign n_25640 =  x_1523 &  n_25639;
assign n_25641 = ~x_1523 & ~n_25639;
assign n_25642 = ~n_25640 & ~n_25641;
assign n_25643 = ~n_25572 & ~n_25573;
assign n_25644 =  x_1524 &  n_25643;
assign n_25645 = ~x_1524 & ~n_25643;
assign n_25646 = ~n_25644 & ~n_25645;
assign n_25647 = ~n_25568 & ~n_25569;
assign n_25648 =  x_1525 &  n_25647;
assign n_25649 = ~x_1525 & ~n_25647;
assign n_25650 = ~n_25648 & ~n_25649;
assign n_25651 = ~n_25564 & ~n_25565;
assign n_25652 =  x_1526 &  n_25651;
assign n_25653 = ~x_1526 & ~n_25651;
assign n_25654 = ~n_25652 & ~n_25653;
assign n_25655 = ~n_25560 & ~n_25561;
assign n_25656 =  x_1527 &  n_25655;
assign n_25657 = ~x_1527 & ~n_25655;
assign n_25658 = ~n_25656 & ~n_25657;
assign n_25659 = ~n_25556 & ~n_25557;
assign n_25660 =  x_1528 &  n_25659;
assign n_25661 = ~x_1528 & ~n_25659;
assign n_25662 = ~n_25660 & ~n_25661;
assign n_25663 = ~n_25552 & ~n_25553;
assign n_25664 =  x_1529 &  n_25663;
assign n_25665 = ~x_1529 & ~n_25663;
assign n_25666 = ~n_25664 & ~n_25665;
assign n_25667 = ~n_25548 & ~n_25549;
assign n_25668 =  x_1530 &  n_25667;
assign n_25669 = ~x_1530 & ~n_25667;
assign n_25670 = ~n_25668 & ~n_25669;
assign n_25671 = ~n_25544 & ~n_25545;
assign n_25672 =  x_1531 &  n_25671;
assign n_25673 = ~x_1531 & ~n_25671;
assign n_25674 = ~n_25672 & ~n_25673;
assign n_25675 = ~n_25540 & ~n_25541;
assign n_25676 =  x_1532 &  n_25675;
assign n_25677 = ~x_1532 & ~n_25675;
assign n_25678 = ~n_25676 & ~n_25677;
assign n_25679 = ~n_25536 & ~n_25537;
assign n_25680 =  x_1533 &  n_25679;
assign n_25681 = ~x_1533 & ~n_25679;
assign n_25682 = ~n_25680 & ~n_25681;
assign n_25683 = ~n_25532 & ~n_25533;
assign n_25684 =  x_1534 &  n_25683;
assign n_25685 = ~x_1534 & ~n_25683;
assign n_25686 = ~n_25684 & ~n_25685;
assign n_25687 = ~n_25528 & ~n_25529;
assign n_25688 =  x_1535 &  n_25687;
assign n_25689 = ~x_1535 & ~n_25687;
assign n_25690 = ~n_25688 & ~n_25689;
assign n_25691 = ~n_25524 & ~n_25525;
assign n_25692 =  x_1536 &  n_25691;
assign n_25693 = ~x_1536 & ~n_25691;
assign n_25694 = ~n_25692 & ~n_25693;
assign n_25695 = ~n_25520 & ~n_25521;
assign n_25696 =  x_1537 &  n_25695;
assign n_25697 = ~x_1537 & ~n_25695;
assign n_25698 = ~n_25696 & ~n_25697;
assign n_25699 = ~n_25516 & ~n_25517;
assign n_25700 =  x_1538 &  n_25699;
assign n_25701 = ~x_1538 & ~n_25699;
assign n_25702 = ~n_25700 & ~n_25701;
assign n_25703 = ~n_25512 & ~n_25513;
assign n_25704 =  x_1539 &  n_25703;
assign n_25705 = ~x_1539 & ~n_25703;
assign n_25706 = ~n_25704 & ~n_25705;
assign n_25707 = ~n_25508 & ~n_25509;
assign n_25708 =  x_1540 &  n_25707;
assign n_25709 = ~x_1540 & ~n_25707;
assign n_25710 = ~n_25708 & ~n_25709;
assign n_25711 = ~n_25504 & ~n_25505;
assign n_25712 =  x_1541 &  n_25711;
assign n_25713 = ~x_1541 & ~n_25711;
assign n_25714 = ~n_25712 & ~n_25713;
assign n_25715 = ~n_25500 & ~n_25501;
assign n_25716 =  x_1542 &  n_25715;
assign n_25717 = ~x_1542 & ~n_25715;
assign n_25718 = ~n_25716 & ~n_25717;
assign n_25719 = ~n_25494 & ~n_25495;
assign n_25720 =  x_1543 &  n_25719;
assign n_25721 = ~x_1543 & ~n_25719;
assign n_25722 = ~n_25720 & ~n_25721;
assign n_25723 = ~n_25487 & ~n_25488;
assign n_25724 = ~n_25491 & ~n_25723;
assign n_25725 = ~n_25487 &  n_25492;
assign n_25726 = ~n_25482 & ~n_25484;
assign n_25727 = ~x_1546 &  x_1610;
assign n_25728 = ~n_25483 & ~n_25727;
assign n_25729 = ~n_25726 &  n_25728;
assign n_25730 = ~n_25725 &  n_25729;
assign n_25731 = ~n_25724 &  n_25730;
assign n_25732 = ~n_25722 &  n_25731;
assign n_25733 = ~n_25718 &  n_25732;
assign n_25734 = ~n_25714 &  n_25733;
assign n_25735 = ~n_25710 &  n_25734;
assign n_25736 = ~n_25706 &  n_25735;
assign n_25737 = ~n_25702 &  n_25736;
assign n_25738 = ~n_25698 &  n_25737;
assign n_25739 = ~n_25694 &  n_25738;
assign n_25740 = ~n_25690 &  n_25739;
assign n_25741 = ~n_25686 &  n_25740;
assign n_25742 = ~n_25682 &  n_25741;
assign n_25743 = ~n_25678 &  n_25742;
assign n_25744 = ~n_25674 &  n_25743;
assign n_25745 = ~n_25670 &  n_25744;
assign n_25746 = ~n_25666 &  n_25745;
assign n_25747 = ~n_25662 &  n_25746;
assign n_25748 = ~n_25658 &  n_25747;
assign n_25749 = ~n_25654 &  n_25748;
assign n_25750 = ~n_25650 &  n_25749;
assign n_25751 = ~n_25646 &  n_25750;
assign n_25752 = ~n_25642 &  n_25751;
assign n_25753 = ~n_25638 &  n_25752;
assign n_25754 = ~n_25634 &  n_25753;
assign n_25755 = ~n_25630 &  n_25754;
assign n_25756 = ~n_25626 &  n_25755;
assign n_25757 = ~n_25622 &  n_25756;
assign n_25758 = ~n_25618 &  n_25757;
assign n_25759 = ~n_25614 &  n_25758;
assign n_25760 = ~n_25609 &  n_25759;
assign n_25761 =  x_1579 &  n_25401;
assign n_25762 = ~n_25610 & ~n_25761;
assign n_25763 = ~n_25400 &  n_25762;
assign n_25764 =  n_25400 & ~n_25762;
assign n_25765 = ~n_25763 & ~n_25764;
assign n_25766 =  n_25613 &  n_25765;
assign n_25767 = ~n_25613 & ~n_25765;
assign n_25768 = ~n_25766 & ~n_25767;
assign n_25769 =  x_1515 & ~n_25768;
assign n_25770 = ~x_1515 &  n_25768;
assign n_25771 = ~n_25769 & ~n_25770;
assign n_25772 =  n_25760 &  n_25771;
assign n_25773 =  n_25320 &  n_25772;
assign n_25774 =  n_13012 &  n_2886;
assign n_25775 =  n_2296 &  n_25774;
assign n_25776 =  n_186 &  n_23891;
assign n_25777 = ~x_2536 & ~x_2537;
assign n_25778 = ~x_2535 &  n_25777;
assign n_25779 = ~x_2534 &  n_25778;
assign n_25780 = ~x_2533 & ~x_2538;
assign n_25781 =  n_25779 &  n_25780;
assign n_25782 = ~x_2532 &  n_25781;
assign n_25783 = ~x_2531 &  n_25782;
assign n_25784 = ~x_2530 &  n_25783;
assign n_25785 = ~x_2529 &  n_25784;
assign n_25786 = ~x_2528 &  n_25785;
assign n_25787 = ~x_2527 &  n_25786;
assign n_25788 = ~x_2526 &  n_25787;
assign n_25789 = ~x_2525 &  n_25788;
assign n_25790 = ~x_2524 &  n_25789;
assign n_25791 = ~x_2523 &  n_25790;
assign n_25792 = ~x_2522 &  n_25791;
assign n_25793 = ~x_2521 &  n_25792;
assign n_25794 = ~x_2520 &  n_25793;
assign n_25795 = ~x_2519 &  n_25794;
assign n_25796 = ~x_2518 &  n_25795;
assign n_25797 = ~x_2517 &  n_25796;
assign n_25798 = ~x_2516 &  n_25797;
assign n_25799 = ~x_2515 &  n_25798;
assign n_25800 = ~x_2514 &  n_25799;
assign n_25801 = ~x_2513 &  n_25800;
assign n_25802 = ~x_2512 &  n_25801;
assign n_25803 = ~x_2511 &  n_25802;
assign n_25804 = ~x_2510 &  n_25803;
assign n_25805 = ~x_2509 &  n_25804;
assign n_25806 =  x_2509 & ~n_25804;
assign n_25807 = ~n_25805 & ~n_25806;
assign n_25808 =  x_2511 & ~n_25802;
assign n_25809 = ~n_25803 & ~n_25808;
assign n_25810 =  x_2513 & ~n_25800;
assign n_25811 = ~n_25801 & ~n_25810;
assign n_25812 =  x_2515 & ~n_25798;
assign n_25813 = ~n_25799 & ~n_25812;
assign n_25814 =  x_2517 & ~n_25796;
assign n_25815 = ~n_25797 & ~n_25814;
assign n_25816 =  x_2519 & ~n_25794;
assign n_25817 = ~n_25795 & ~n_25816;
assign n_25818 =  x_2521 & ~n_25792;
assign n_25819 = ~n_25793 & ~n_25818;
assign n_25820 =  x_2523 & ~n_25790;
assign n_25821 = ~n_25791 & ~n_25820;
assign n_25822 =  x_2525 & ~n_25788;
assign n_25823 = ~n_25789 & ~n_25822;
assign n_25824 =  x_2527 & ~n_25786;
assign n_25825 = ~n_25787 & ~n_25824;
assign n_25826 =  x_2529 & ~n_25784;
assign n_25827 = ~n_25785 & ~n_25826;
assign n_25828 =  x_2531 & ~n_25782;
assign n_25829 = ~n_25783 & ~n_25828;
assign n_25830 = ~x_2533 &  x_2538;
assign n_25831 =  n_25779 &  n_25830;
assign n_25832 = ~x_2532 &  n_25831;
assign n_25833 =  n_25829 &  n_25832;
assign n_25834 = ~x_2530 &  n_25833;
assign n_25835 =  n_25827 &  n_25834;
assign n_25836 = ~x_2528 &  n_25835;
assign n_25837 =  n_25825 &  n_25836;
assign n_25838 = ~x_2526 &  n_25837;
assign n_25839 =  n_25823 &  n_25838;
assign n_25840 = ~x_2524 &  n_25839;
assign n_25841 =  n_25821 &  n_25840;
assign n_25842 = ~x_2522 &  n_25841;
assign n_25843 =  n_25819 &  n_25842;
assign n_25844 = ~x_2520 &  n_25843;
assign n_25845 =  n_25817 &  n_25844;
assign n_25846 = ~x_2518 &  n_25845;
assign n_25847 =  n_25815 &  n_25846;
assign n_25848 = ~x_2516 &  n_25847;
assign n_25849 =  n_25813 &  n_25848;
assign n_25850 = ~x_2514 &  n_25849;
assign n_25851 =  n_25811 &  n_25850;
assign n_25852 = ~x_2512 &  n_25851;
assign n_25853 =  n_25809 &  n_25852;
assign n_25854 = ~x_2510 &  n_25853;
assign n_25855 =  n_25807 &  n_25854;
assign n_25856 = ~x_2508 &  n_25855;
assign n_25857 = ~x_2508 &  n_25805;
assign n_25858 =  x_2508 & ~n_25805;
assign n_25859 = ~n_25857 & ~n_25858;
assign n_25860 = ~n_25855 & ~n_25859;
assign n_25861 = ~n_25856 & ~n_25860;
assign n_25862 = ~n_25807 & ~n_25854;
assign n_25863 = ~n_25855 & ~n_25862;
assign n_25864 =  x_2510 & ~n_25803;
assign n_25865 = ~n_25804 & ~n_25864;
assign n_25866 = ~n_25853 & ~n_25865;
assign n_25867 = ~n_25854 & ~n_25866;
assign n_25868 = ~n_25809 & ~n_25852;
assign n_25869 = ~n_25853 & ~n_25868;
assign n_25870 =  x_2512 & ~n_25801;
assign n_25871 = ~n_25802 & ~n_25870;
assign n_25872 = ~n_25851 & ~n_25871;
assign n_25873 = ~n_25852 & ~n_25872;
assign n_25874 = ~n_25811 & ~n_25850;
assign n_25875 = ~n_25851 & ~n_25874;
assign n_25876 =  x_2514 & ~n_25799;
assign n_25877 = ~n_25800 & ~n_25876;
assign n_25878 = ~n_25849 & ~n_25877;
assign n_25879 = ~n_25850 & ~n_25878;
assign n_25880 = ~n_25813 & ~n_25848;
assign n_25881 = ~n_25849 & ~n_25880;
assign n_25882 =  x_2516 & ~n_25797;
assign n_25883 = ~n_25798 & ~n_25882;
assign n_25884 = ~n_25847 & ~n_25883;
assign n_25885 = ~n_25848 & ~n_25884;
assign n_25886 = ~n_25815 & ~n_25846;
assign n_25887 = ~n_25847 & ~n_25886;
assign n_25888 =  x_2518 & ~n_25795;
assign n_25889 = ~n_25796 & ~n_25888;
assign n_25890 = ~n_25845 & ~n_25889;
assign n_25891 = ~n_25846 & ~n_25890;
assign n_25892 = ~n_25817 & ~n_25844;
assign n_25893 = ~n_25845 & ~n_25892;
assign n_25894 =  x_2520 & ~n_25793;
assign n_25895 = ~n_25794 & ~n_25894;
assign n_25896 = ~n_25843 & ~n_25895;
assign n_25897 = ~n_25844 & ~n_25896;
assign n_25898 = ~n_25819 & ~n_25842;
assign n_25899 = ~n_25843 & ~n_25898;
assign n_25900 =  x_2522 & ~n_25791;
assign n_25901 = ~n_25792 & ~n_25900;
assign n_25902 = ~n_25841 & ~n_25901;
assign n_25903 = ~n_25842 & ~n_25902;
assign n_25904 = ~n_25821 & ~n_25840;
assign n_25905 = ~n_25841 & ~n_25904;
assign n_25906 =  x_2524 & ~n_25789;
assign n_25907 = ~n_25790 & ~n_25906;
assign n_25908 = ~n_25839 & ~n_25907;
assign n_25909 = ~n_25840 & ~n_25908;
assign n_25910 = ~n_25823 & ~n_25838;
assign n_25911 = ~n_25839 & ~n_25910;
assign n_25912 =  x_2526 & ~n_25787;
assign n_25913 = ~n_25788 & ~n_25912;
assign n_25914 = ~n_25837 & ~n_25913;
assign n_25915 = ~n_25838 & ~n_25914;
assign n_25916 = ~n_25825 & ~n_25836;
assign n_25917 = ~n_25837 & ~n_25916;
assign n_25918 =  x_2528 & ~n_25785;
assign n_25919 = ~n_25786 & ~n_25918;
assign n_25920 = ~n_25835 & ~n_25919;
assign n_25921 = ~n_25836 & ~n_25920;
assign n_25922 = ~n_25827 & ~n_25834;
assign n_25923 = ~n_25835 & ~n_25922;
assign n_25924 =  x_2530 & ~n_25783;
assign n_25925 = ~n_25784 & ~n_25924;
assign n_25926 = ~n_25833 & ~n_25925;
assign n_25927 = ~n_25834 & ~n_25926;
assign n_25928 = ~n_25829 & ~n_25832;
assign n_25929 = ~n_25833 & ~n_25928;
assign n_25930 = ~n_25781 & ~n_25831;
assign n_25931 =  x_2532 & ~n_25930;
assign n_25932 = ~x_2532 &  n_25930;
assign n_25933 = ~n_25931 & ~n_25932;
assign n_25934 =  x_2533 & ~n_25779;
assign n_25935 =  n_25930 & ~n_25934;
assign n_25936 =  x_2535 & ~n_25777;
assign n_25937 = ~n_25778 & ~n_25936;
assign n_25938 = ~x_2505 & ~x_2537;
assign n_25939 =  x_2506 & ~x_2538;
assign n_25940 =  x_2505 &  x_2537;
assign n_25941 = ~n_25939 & ~n_25940;
assign n_25942 = ~n_25938 & ~n_25941;
assign n_25943 = ~x_2504 & ~n_25942;
assign n_25944 =  x_2536 & ~x_2537;
assign n_25945 = ~x_2536 &  x_2537;
assign n_25946 = ~n_25944 & ~n_25945;
assign n_25947 =  x_2504 &  n_25942;
assign n_25948 =  n_25946 & ~n_25947;
assign n_25949 = ~n_25943 & ~n_25948;
assign n_25950 = ~n_25937 & ~n_25949;
assign n_25951 =  n_25937 &  n_25949;
assign n_25952 = ~x_2503 & ~n_25951;
assign n_25953 = ~n_25950 & ~n_25952;
assign n_25954 =  x_2534 & ~n_25778;
assign n_25955 = ~n_25779 & ~n_25954;
assign n_25956 = ~n_25953 & ~n_25955;
assign n_25957 =  n_25953 &  n_25955;
assign n_25958 = ~x_2502 & ~n_25957;
assign n_25959 = ~n_25956 & ~n_25958;
assign n_25960 = ~n_25935 & ~n_25959;
assign n_25961 =  n_25935 &  n_25959;
assign n_25962 = ~x_2501 & ~n_25961;
assign n_25963 = ~n_25960 & ~n_25962;
assign n_25964 =  n_25933 & ~n_25963;
assign n_25965 = ~n_25933 &  n_25963;
assign n_25966 = ~x_2500 & ~n_25965;
assign n_25967 = ~n_25964 & ~n_25966;
assign n_25968 = ~n_25929 & ~n_25967;
assign n_25969 =  n_25929 &  n_25967;
assign n_25970 = ~x_2499 & ~n_25969;
assign n_25971 = ~n_25968 & ~n_25970;
assign n_25972 = ~n_25927 & ~n_25971;
assign n_25973 =  n_25927 &  n_25971;
assign n_25974 = ~x_2498 & ~n_25973;
assign n_25975 = ~n_25972 & ~n_25974;
assign n_25976 = ~n_25923 & ~n_25975;
assign n_25977 =  n_25923 &  n_25975;
assign n_25978 = ~x_2497 & ~n_25977;
assign n_25979 = ~n_25976 & ~n_25978;
assign n_25980 = ~n_25921 & ~n_25979;
assign n_25981 =  n_25921 &  n_25979;
assign n_25982 = ~x_2496 & ~n_25981;
assign n_25983 = ~n_25980 & ~n_25982;
assign n_25984 = ~n_25917 & ~n_25983;
assign n_25985 =  n_25917 &  n_25983;
assign n_25986 = ~x_2495 & ~n_25985;
assign n_25987 = ~n_25984 & ~n_25986;
assign n_25988 = ~n_25915 & ~n_25987;
assign n_25989 =  n_25915 &  n_25987;
assign n_25990 = ~x_2494 & ~n_25989;
assign n_25991 = ~n_25988 & ~n_25990;
assign n_25992 = ~n_25911 & ~n_25991;
assign n_25993 =  n_25911 &  n_25991;
assign n_25994 = ~x_2493 & ~n_25993;
assign n_25995 = ~n_25992 & ~n_25994;
assign n_25996 = ~n_25909 & ~n_25995;
assign n_25997 =  n_25909 &  n_25995;
assign n_25998 = ~x_2492 & ~n_25997;
assign n_25999 = ~n_25996 & ~n_25998;
assign n_26000 = ~n_25905 & ~n_25999;
assign n_26001 =  n_25905 &  n_25999;
assign n_26002 = ~x_2491 & ~n_26001;
assign n_26003 = ~n_26000 & ~n_26002;
assign n_26004 = ~n_25903 & ~n_26003;
assign n_26005 =  n_25903 &  n_26003;
assign n_26006 = ~x_2490 & ~n_26005;
assign n_26007 = ~n_26004 & ~n_26006;
assign n_26008 = ~n_25899 & ~n_26007;
assign n_26009 =  n_25899 &  n_26007;
assign n_26010 = ~x_2489 & ~n_26009;
assign n_26011 = ~n_26008 & ~n_26010;
assign n_26012 = ~n_25897 & ~n_26011;
assign n_26013 =  n_25897 &  n_26011;
assign n_26014 = ~x_2488 & ~n_26013;
assign n_26015 = ~n_26012 & ~n_26014;
assign n_26016 = ~n_25893 & ~n_26015;
assign n_26017 =  n_25893 &  n_26015;
assign n_26018 = ~x_2487 & ~n_26017;
assign n_26019 = ~n_26016 & ~n_26018;
assign n_26020 = ~n_25891 & ~n_26019;
assign n_26021 =  n_25891 &  n_26019;
assign n_26022 = ~x_2486 & ~n_26021;
assign n_26023 = ~n_26020 & ~n_26022;
assign n_26024 = ~n_25887 & ~n_26023;
assign n_26025 =  n_25887 &  n_26023;
assign n_26026 = ~x_2485 & ~n_26025;
assign n_26027 = ~n_26024 & ~n_26026;
assign n_26028 = ~n_25885 & ~n_26027;
assign n_26029 =  n_25885 &  n_26027;
assign n_26030 = ~x_2484 & ~n_26029;
assign n_26031 = ~n_26028 & ~n_26030;
assign n_26032 = ~n_25881 & ~n_26031;
assign n_26033 =  n_25881 &  n_26031;
assign n_26034 = ~x_2483 & ~n_26033;
assign n_26035 = ~n_26032 & ~n_26034;
assign n_26036 = ~n_25879 & ~n_26035;
assign n_26037 =  n_25879 &  n_26035;
assign n_26038 = ~x_2482 & ~n_26037;
assign n_26039 = ~n_26036 & ~n_26038;
assign n_26040 = ~n_25875 & ~n_26039;
assign n_26041 =  n_25875 &  n_26039;
assign n_26042 = ~x_2481 & ~n_26041;
assign n_26043 = ~n_26040 & ~n_26042;
assign n_26044 = ~n_25873 & ~n_26043;
assign n_26045 =  n_25873 &  n_26043;
assign n_26046 = ~x_2480 & ~n_26045;
assign n_26047 = ~n_26044 & ~n_26046;
assign n_26048 = ~n_25869 & ~n_26047;
assign n_26049 =  n_25869 &  n_26047;
assign n_26050 = ~x_2479 & ~n_26049;
assign n_26051 = ~n_26048 & ~n_26050;
assign n_26052 = ~n_25867 & ~n_26051;
assign n_26053 =  n_25867 &  n_26051;
assign n_26054 = ~x_2478 & ~n_26053;
assign n_26055 = ~n_26052 & ~n_26054;
assign n_26056 = ~n_25863 & ~n_26055;
assign n_26057 =  n_25863 &  n_26055;
assign n_26058 = ~x_2477 & ~n_26057;
assign n_26059 = ~n_26056 & ~n_26058;
assign n_26060 = ~n_25861 & ~n_26059;
assign n_26061 =  n_25861 &  n_26059;
assign n_26062 = ~n_26060 & ~n_26061;
assign n_26063 = ~x_2476 & ~n_26062;
assign n_26064 =  x_2476 &  n_26062;
assign n_26065 = ~n_26063 & ~n_26064;
assign n_26066 = ~n_26056 & ~n_26057;
assign n_26067 =  x_2477 &  n_26066;
assign n_26068 = ~x_2477 & ~n_26066;
assign n_26069 = ~n_26067 & ~n_26068;
assign n_26070 = ~n_26052 & ~n_26053;
assign n_26071 =  x_2478 &  n_26070;
assign n_26072 = ~x_2478 & ~n_26070;
assign n_26073 = ~n_26071 & ~n_26072;
assign n_26074 = ~n_26048 & ~n_26049;
assign n_26075 =  x_2479 &  n_26074;
assign n_26076 = ~x_2479 & ~n_26074;
assign n_26077 = ~n_26075 & ~n_26076;
assign n_26078 = ~n_26044 & ~n_26045;
assign n_26079 =  x_2480 &  n_26078;
assign n_26080 = ~x_2480 & ~n_26078;
assign n_26081 = ~n_26079 & ~n_26080;
assign n_26082 = ~n_26040 & ~n_26041;
assign n_26083 =  x_2481 &  n_26082;
assign n_26084 = ~x_2481 & ~n_26082;
assign n_26085 = ~n_26083 & ~n_26084;
assign n_26086 = ~n_26036 & ~n_26037;
assign n_26087 =  x_2482 &  n_26086;
assign n_26088 = ~x_2482 & ~n_26086;
assign n_26089 = ~n_26087 & ~n_26088;
assign n_26090 = ~n_26032 & ~n_26033;
assign n_26091 =  x_2483 &  n_26090;
assign n_26092 = ~x_2483 & ~n_26090;
assign n_26093 = ~n_26091 & ~n_26092;
assign n_26094 = ~n_26028 & ~n_26029;
assign n_26095 =  x_2484 &  n_26094;
assign n_26096 = ~x_2484 & ~n_26094;
assign n_26097 = ~n_26095 & ~n_26096;
assign n_26098 = ~n_26024 & ~n_26025;
assign n_26099 =  x_2485 &  n_26098;
assign n_26100 = ~x_2485 & ~n_26098;
assign n_26101 = ~n_26099 & ~n_26100;
assign n_26102 = ~n_26020 & ~n_26021;
assign n_26103 =  x_2486 &  n_26102;
assign n_26104 = ~x_2486 & ~n_26102;
assign n_26105 = ~n_26103 & ~n_26104;
assign n_26106 = ~n_26016 & ~n_26017;
assign n_26107 =  x_2487 &  n_26106;
assign n_26108 = ~x_2487 & ~n_26106;
assign n_26109 = ~n_26107 & ~n_26108;
assign n_26110 = ~n_26012 & ~n_26013;
assign n_26111 =  x_2488 &  n_26110;
assign n_26112 = ~x_2488 & ~n_26110;
assign n_26113 = ~n_26111 & ~n_26112;
assign n_26114 = ~n_26008 & ~n_26009;
assign n_26115 =  x_2489 &  n_26114;
assign n_26116 = ~x_2489 & ~n_26114;
assign n_26117 = ~n_26115 & ~n_26116;
assign n_26118 = ~n_26004 & ~n_26005;
assign n_26119 =  x_2490 &  n_26118;
assign n_26120 = ~x_2490 & ~n_26118;
assign n_26121 = ~n_26119 & ~n_26120;
assign n_26122 = ~n_26000 & ~n_26001;
assign n_26123 =  x_2491 &  n_26122;
assign n_26124 = ~x_2491 & ~n_26122;
assign n_26125 = ~n_26123 & ~n_26124;
assign n_26126 = ~n_25996 & ~n_25997;
assign n_26127 =  x_2492 &  n_26126;
assign n_26128 = ~x_2492 & ~n_26126;
assign n_26129 = ~n_26127 & ~n_26128;
assign n_26130 = ~n_25992 & ~n_25993;
assign n_26131 =  x_2493 &  n_26130;
assign n_26132 = ~x_2493 & ~n_26130;
assign n_26133 = ~n_26131 & ~n_26132;
assign n_26134 = ~n_25988 & ~n_25989;
assign n_26135 =  x_2494 &  n_26134;
assign n_26136 = ~x_2494 & ~n_26134;
assign n_26137 = ~n_26135 & ~n_26136;
assign n_26138 = ~n_25984 & ~n_25985;
assign n_26139 =  x_2495 &  n_26138;
assign n_26140 = ~x_2495 & ~n_26138;
assign n_26141 = ~n_26139 & ~n_26140;
assign n_26142 = ~n_25980 & ~n_25981;
assign n_26143 =  x_2496 &  n_26142;
assign n_26144 = ~x_2496 & ~n_26142;
assign n_26145 = ~n_26143 & ~n_26144;
assign n_26146 = ~n_25976 & ~n_25977;
assign n_26147 =  x_2497 &  n_26146;
assign n_26148 = ~x_2497 & ~n_26146;
assign n_26149 = ~n_26147 & ~n_26148;
assign n_26150 = ~n_25972 & ~n_25973;
assign n_26151 =  x_2498 &  n_26150;
assign n_26152 = ~x_2498 & ~n_26150;
assign n_26153 = ~n_26151 & ~n_26152;
assign n_26154 = ~n_25968 & ~n_25969;
assign n_26155 =  x_2499 &  n_26154;
assign n_26156 = ~x_2499 & ~n_26154;
assign n_26157 = ~n_26155 & ~n_26156;
assign n_26158 = ~n_25964 & ~n_25965;
assign n_26159 =  x_2500 &  n_26158;
assign n_26160 = ~x_2500 & ~n_26158;
assign n_26161 = ~n_26159 & ~n_26160;
assign n_26162 = ~n_25960 & ~n_25961;
assign n_26163 =  x_2501 &  n_26162;
assign n_26164 = ~x_2501 & ~n_26162;
assign n_26165 = ~n_26163 & ~n_26164;
assign n_26166 = ~n_25956 & ~n_25957;
assign n_26167 =  x_2502 &  n_26166;
assign n_26168 = ~x_2502 & ~n_26166;
assign n_26169 = ~n_26167 & ~n_26168;
assign n_26170 = ~n_25950 & ~n_25951;
assign n_26171 =  x_2503 &  n_26170;
assign n_26172 = ~x_2503 & ~n_26170;
assign n_26173 = ~n_26171 & ~n_26172;
assign n_26174 = ~n_25943 & ~n_25947;
assign n_26175 = ~n_25946 & ~n_26174;
assign n_26176 = ~n_25943 &  n_25948;
assign n_26177 = ~n_25938 & ~n_25940;
assign n_26178 = ~x_2506 &  x_2538;
assign n_26179 = ~n_25939 & ~n_26178;
assign n_26180 = ~n_26177 &  n_26179;
assign n_26181 = ~n_26176 &  n_26180;
assign n_26182 = ~n_26175 &  n_26181;
assign n_26183 = ~n_26173 &  n_26182;
assign n_26184 = ~n_26169 &  n_26183;
assign n_26185 = ~n_26165 &  n_26184;
assign n_26186 = ~n_26161 &  n_26185;
assign n_26187 = ~n_26157 &  n_26186;
assign n_26188 = ~n_26153 &  n_26187;
assign n_26189 = ~n_26149 &  n_26188;
assign n_26190 = ~n_26145 &  n_26189;
assign n_26191 = ~n_26141 &  n_26190;
assign n_26192 = ~n_26137 &  n_26191;
assign n_26193 = ~n_26133 &  n_26192;
assign n_26194 = ~n_26129 &  n_26193;
assign n_26195 = ~n_26125 &  n_26194;
assign n_26196 = ~n_26121 &  n_26195;
assign n_26197 = ~n_26117 &  n_26196;
assign n_26198 = ~n_26113 &  n_26197;
assign n_26199 = ~n_26109 &  n_26198;
assign n_26200 = ~n_26105 &  n_26199;
assign n_26201 = ~n_26101 &  n_26200;
assign n_26202 = ~n_26097 &  n_26201;
assign n_26203 = ~n_26093 &  n_26202;
assign n_26204 = ~n_26089 &  n_26203;
assign n_26205 = ~n_26085 &  n_26204;
assign n_26206 = ~n_26081 &  n_26205;
assign n_26207 = ~n_26077 &  n_26206;
assign n_26208 = ~n_26073 &  n_26207;
assign n_26209 = ~n_26069 &  n_26208;
assign n_26210 = ~n_26065 &  n_26209;
assign n_26211 = ~x_2507 & ~n_25857;
assign n_26212 =  x_2507 &  n_25857;
assign n_26213 = ~n_26211 & ~n_26212;
assign n_26214 = ~n_25856 &  n_26213;
assign n_26215 =  n_25856 & ~n_26213;
assign n_26216 = ~n_26214 & ~n_26215;
assign n_26217 = ~x_2476 & ~n_26061;
assign n_26218 = ~n_26060 & ~n_26217;
assign n_26219 =  n_26216 &  n_26218;
assign n_26220 = ~n_26216 & ~n_26218;
assign n_26221 = ~n_26219 & ~n_26220;
assign n_26222 =  x_2475 & ~n_26221;
assign n_26223 = ~x_2475 &  n_26221;
assign n_26224 = ~n_26222 & ~n_26223;
assign n_26225 =  n_26210 &  n_26224;
assign n_26226 =  n_25776 &  n_26225;
assign n_26227 = ~n_25775 & ~n_26226;
assign n_26228 = ~n_25773 &  n_26227;
assign n_26229 =  n_980 &  n_12226;
assign n_26230 = ~x_1288 & ~x_1289;
assign n_26231 = ~x_1287 &  n_26230;
assign n_26232 = ~x_1286 &  n_26231;
assign n_26233 = ~x_1285 & ~x_1290;
assign n_26234 =  n_26232 &  n_26233;
assign n_26235 = ~x_1284 &  n_26234;
assign n_26236 = ~x_1283 &  n_26235;
assign n_26237 = ~x_1282 &  n_26236;
assign n_26238 = ~x_1281 &  n_26237;
assign n_26239 = ~x_1280 &  n_26238;
assign n_26240 = ~x_1279 &  n_26239;
assign n_26241 = ~x_1278 &  n_26240;
assign n_26242 = ~x_1277 &  n_26241;
assign n_26243 = ~x_1276 &  n_26242;
assign n_26244 = ~x_1275 &  n_26243;
assign n_26245 = ~x_1274 &  n_26244;
assign n_26246 = ~x_1273 &  n_26245;
assign n_26247 = ~x_1272 &  n_26246;
assign n_26248 = ~x_1271 &  n_26247;
assign n_26249 = ~x_1270 &  n_26248;
assign n_26250 = ~x_1269 &  n_26249;
assign n_26251 = ~x_1268 &  n_26250;
assign n_26252 = ~x_1267 &  n_26251;
assign n_26253 = ~x_1266 &  n_26252;
assign n_26254 = ~x_1265 &  n_26253;
assign n_26255 = ~x_1264 &  n_26254;
assign n_26256 = ~x_1263 &  n_26255;
assign n_26257 = ~x_1262 &  n_26256;
assign n_26258 = ~x_1261 &  n_26257;
assign n_26259 =  x_1261 & ~n_26257;
assign n_26260 = ~n_26258 & ~n_26259;
assign n_26261 =  x_1263 & ~n_26255;
assign n_26262 = ~n_26256 & ~n_26261;
assign n_26263 =  x_1265 & ~n_26253;
assign n_26264 = ~n_26254 & ~n_26263;
assign n_26265 =  x_1267 & ~n_26251;
assign n_26266 = ~n_26252 & ~n_26265;
assign n_26267 =  x_1269 & ~n_26249;
assign n_26268 = ~n_26250 & ~n_26267;
assign n_26269 =  x_1271 & ~n_26247;
assign n_26270 = ~n_26248 & ~n_26269;
assign n_26271 =  x_1273 & ~n_26245;
assign n_26272 = ~n_26246 & ~n_26271;
assign n_26273 =  x_1275 & ~n_26243;
assign n_26274 = ~n_26244 & ~n_26273;
assign n_26275 =  x_1277 & ~n_26241;
assign n_26276 = ~n_26242 & ~n_26275;
assign n_26277 =  x_1279 & ~n_26239;
assign n_26278 = ~n_26240 & ~n_26277;
assign n_26279 =  x_1281 & ~n_26237;
assign n_26280 = ~n_26238 & ~n_26279;
assign n_26281 =  x_1283 & ~n_26235;
assign n_26282 = ~n_26236 & ~n_26281;
assign n_26283 = ~x_1285 &  x_1290;
assign n_26284 =  n_26232 &  n_26283;
assign n_26285 = ~x_1284 &  n_26284;
assign n_26286 =  n_26282 &  n_26285;
assign n_26287 = ~x_1282 &  n_26286;
assign n_26288 =  n_26280 &  n_26287;
assign n_26289 = ~x_1280 &  n_26288;
assign n_26290 =  n_26278 &  n_26289;
assign n_26291 = ~x_1278 &  n_26290;
assign n_26292 =  n_26276 &  n_26291;
assign n_26293 = ~x_1276 &  n_26292;
assign n_26294 =  n_26274 &  n_26293;
assign n_26295 = ~x_1274 &  n_26294;
assign n_26296 =  n_26272 &  n_26295;
assign n_26297 = ~x_1272 &  n_26296;
assign n_26298 =  n_26270 &  n_26297;
assign n_26299 = ~x_1270 &  n_26298;
assign n_26300 =  n_26268 &  n_26299;
assign n_26301 = ~x_1268 &  n_26300;
assign n_26302 =  n_26266 &  n_26301;
assign n_26303 = ~x_1266 &  n_26302;
assign n_26304 =  n_26264 &  n_26303;
assign n_26305 = ~x_1264 &  n_26304;
assign n_26306 =  n_26262 &  n_26305;
assign n_26307 = ~x_1262 &  n_26306;
assign n_26308 =  n_26260 &  n_26307;
assign n_26309 = ~x_1260 &  n_26308;
assign n_26310 = ~x_1260 &  n_26258;
assign n_26311 =  x_1260 & ~n_26258;
assign n_26312 = ~n_26310 & ~n_26311;
assign n_26313 = ~n_26308 & ~n_26312;
assign n_26314 = ~n_26309 & ~n_26313;
assign n_26315 = ~n_26260 & ~n_26307;
assign n_26316 = ~n_26308 & ~n_26315;
assign n_26317 =  x_1262 & ~n_26256;
assign n_26318 = ~n_26257 & ~n_26317;
assign n_26319 = ~n_26306 & ~n_26318;
assign n_26320 = ~n_26307 & ~n_26319;
assign n_26321 = ~n_26262 & ~n_26305;
assign n_26322 = ~n_26306 & ~n_26321;
assign n_26323 =  x_1264 & ~n_26254;
assign n_26324 = ~n_26255 & ~n_26323;
assign n_26325 = ~n_26304 & ~n_26324;
assign n_26326 = ~n_26305 & ~n_26325;
assign n_26327 = ~n_26264 & ~n_26303;
assign n_26328 = ~n_26304 & ~n_26327;
assign n_26329 =  x_1266 & ~n_26252;
assign n_26330 = ~n_26253 & ~n_26329;
assign n_26331 = ~n_26302 & ~n_26330;
assign n_26332 = ~n_26303 & ~n_26331;
assign n_26333 = ~n_26266 & ~n_26301;
assign n_26334 = ~n_26302 & ~n_26333;
assign n_26335 =  x_1268 & ~n_26250;
assign n_26336 = ~n_26251 & ~n_26335;
assign n_26337 = ~n_26300 & ~n_26336;
assign n_26338 = ~n_26301 & ~n_26337;
assign n_26339 = ~n_26268 & ~n_26299;
assign n_26340 = ~n_26300 & ~n_26339;
assign n_26341 =  x_1270 & ~n_26248;
assign n_26342 = ~n_26249 & ~n_26341;
assign n_26343 = ~n_26298 & ~n_26342;
assign n_26344 = ~n_26299 & ~n_26343;
assign n_26345 = ~n_26270 & ~n_26297;
assign n_26346 = ~n_26298 & ~n_26345;
assign n_26347 =  x_1272 & ~n_26246;
assign n_26348 = ~n_26247 & ~n_26347;
assign n_26349 = ~n_26296 & ~n_26348;
assign n_26350 = ~n_26297 & ~n_26349;
assign n_26351 = ~n_26272 & ~n_26295;
assign n_26352 = ~n_26296 & ~n_26351;
assign n_26353 =  x_1274 & ~n_26244;
assign n_26354 = ~n_26245 & ~n_26353;
assign n_26355 = ~n_26294 & ~n_26354;
assign n_26356 = ~n_26295 & ~n_26355;
assign n_26357 = ~n_26274 & ~n_26293;
assign n_26358 = ~n_26294 & ~n_26357;
assign n_26359 =  x_1276 & ~n_26242;
assign n_26360 = ~n_26243 & ~n_26359;
assign n_26361 = ~n_26292 & ~n_26360;
assign n_26362 = ~n_26293 & ~n_26361;
assign n_26363 = ~n_26276 & ~n_26291;
assign n_26364 = ~n_26292 & ~n_26363;
assign n_26365 =  x_1278 & ~n_26240;
assign n_26366 = ~n_26241 & ~n_26365;
assign n_26367 = ~n_26290 & ~n_26366;
assign n_26368 = ~n_26291 & ~n_26367;
assign n_26369 = ~n_26278 & ~n_26289;
assign n_26370 = ~n_26290 & ~n_26369;
assign n_26371 =  x_1280 & ~n_26238;
assign n_26372 = ~n_26239 & ~n_26371;
assign n_26373 = ~n_26288 & ~n_26372;
assign n_26374 = ~n_26289 & ~n_26373;
assign n_26375 = ~n_26280 & ~n_26287;
assign n_26376 = ~n_26288 & ~n_26375;
assign n_26377 =  x_1282 & ~n_26236;
assign n_26378 = ~n_26237 & ~n_26377;
assign n_26379 = ~n_26286 & ~n_26378;
assign n_26380 = ~n_26287 & ~n_26379;
assign n_26381 = ~n_26282 & ~n_26285;
assign n_26382 = ~n_26286 & ~n_26381;
assign n_26383 = ~n_26234 & ~n_26284;
assign n_26384 =  x_1284 & ~n_26383;
assign n_26385 = ~x_1284 &  n_26383;
assign n_26386 = ~n_26384 & ~n_26385;
assign n_26387 =  x_1285 & ~n_26232;
assign n_26388 =  n_26383 & ~n_26387;
assign n_26389 =  x_1287 & ~n_26230;
assign n_26390 = ~n_26231 & ~n_26389;
assign n_26391 = ~x_1257 & ~x_1289;
assign n_26392 =  x_1258 & ~x_1290;
assign n_26393 =  x_1257 &  x_1289;
assign n_26394 = ~n_26392 & ~n_26393;
assign n_26395 = ~n_26391 & ~n_26394;
assign n_26396 = ~x_1256 & ~n_26395;
assign n_26397 =  x_1288 & ~x_1289;
assign n_26398 = ~x_1288 &  x_1289;
assign n_26399 = ~n_26397 & ~n_26398;
assign n_26400 =  x_1256 &  n_26395;
assign n_26401 =  n_26399 & ~n_26400;
assign n_26402 = ~n_26396 & ~n_26401;
assign n_26403 = ~n_26390 & ~n_26402;
assign n_26404 =  n_26390 &  n_26402;
assign n_26405 = ~x_1255 & ~n_26404;
assign n_26406 = ~n_26403 & ~n_26405;
assign n_26407 =  x_1286 & ~n_26231;
assign n_26408 = ~n_26232 & ~n_26407;
assign n_26409 = ~n_26406 & ~n_26408;
assign n_26410 =  n_26406 &  n_26408;
assign n_26411 = ~x_1254 & ~n_26410;
assign n_26412 = ~n_26409 & ~n_26411;
assign n_26413 = ~n_26388 & ~n_26412;
assign n_26414 =  n_26388 &  n_26412;
assign n_26415 = ~x_1253 & ~n_26414;
assign n_26416 = ~n_26413 & ~n_26415;
assign n_26417 =  n_26386 & ~n_26416;
assign n_26418 = ~n_26386 &  n_26416;
assign n_26419 = ~x_1252 & ~n_26418;
assign n_26420 = ~n_26417 & ~n_26419;
assign n_26421 = ~n_26382 & ~n_26420;
assign n_26422 =  n_26382 &  n_26420;
assign n_26423 = ~x_1251 & ~n_26422;
assign n_26424 = ~n_26421 & ~n_26423;
assign n_26425 = ~n_26380 & ~n_26424;
assign n_26426 =  n_26380 &  n_26424;
assign n_26427 = ~x_1250 & ~n_26426;
assign n_26428 = ~n_26425 & ~n_26427;
assign n_26429 = ~n_26376 & ~n_26428;
assign n_26430 =  n_26376 &  n_26428;
assign n_26431 = ~x_1249 & ~n_26430;
assign n_26432 = ~n_26429 & ~n_26431;
assign n_26433 = ~n_26374 & ~n_26432;
assign n_26434 =  n_26374 &  n_26432;
assign n_26435 = ~x_1248 & ~n_26434;
assign n_26436 = ~n_26433 & ~n_26435;
assign n_26437 = ~n_26370 & ~n_26436;
assign n_26438 =  n_26370 &  n_26436;
assign n_26439 = ~x_1247 & ~n_26438;
assign n_26440 = ~n_26437 & ~n_26439;
assign n_26441 = ~n_26368 & ~n_26440;
assign n_26442 =  n_26368 &  n_26440;
assign n_26443 = ~x_1246 & ~n_26442;
assign n_26444 = ~n_26441 & ~n_26443;
assign n_26445 = ~n_26364 & ~n_26444;
assign n_26446 =  n_26364 &  n_26444;
assign n_26447 = ~x_1245 & ~n_26446;
assign n_26448 = ~n_26445 & ~n_26447;
assign n_26449 = ~n_26362 & ~n_26448;
assign n_26450 =  n_26362 &  n_26448;
assign n_26451 = ~x_1244 & ~n_26450;
assign n_26452 = ~n_26449 & ~n_26451;
assign n_26453 = ~n_26358 & ~n_26452;
assign n_26454 =  n_26358 &  n_26452;
assign n_26455 = ~x_1243 & ~n_26454;
assign n_26456 = ~n_26453 & ~n_26455;
assign n_26457 = ~n_26356 & ~n_26456;
assign n_26458 =  n_26356 &  n_26456;
assign n_26459 = ~x_1242 & ~n_26458;
assign n_26460 = ~n_26457 & ~n_26459;
assign n_26461 = ~n_26352 & ~n_26460;
assign n_26462 =  n_26352 &  n_26460;
assign n_26463 = ~x_1241 & ~n_26462;
assign n_26464 = ~n_26461 & ~n_26463;
assign n_26465 = ~n_26350 & ~n_26464;
assign n_26466 =  n_26350 &  n_26464;
assign n_26467 = ~x_1240 & ~n_26466;
assign n_26468 = ~n_26465 & ~n_26467;
assign n_26469 = ~n_26346 & ~n_26468;
assign n_26470 =  n_26346 &  n_26468;
assign n_26471 = ~x_1239 & ~n_26470;
assign n_26472 = ~n_26469 & ~n_26471;
assign n_26473 = ~n_26344 & ~n_26472;
assign n_26474 =  n_26344 &  n_26472;
assign n_26475 = ~x_1238 & ~n_26474;
assign n_26476 = ~n_26473 & ~n_26475;
assign n_26477 = ~n_26340 & ~n_26476;
assign n_26478 =  n_26340 &  n_26476;
assign n_26479 = ~x_1237 & ~n_26478;
assign n_26480 = ~n_26477 & ~n_26479;
assign n_26481 = ~n_26338 & ~n_26480;
assign n_26482 =  n_26338 &  n_26480;
assign n_26483 = ~x_1236 & ~n_26482;
assign n_26484 = ~n_26481 & ~n_26483;
assign n_26485 = ~n_26334 & ~n_26484;
assign n_26486 =  n_26334 &  n_26484;
assign n_26487 = ~x_1235 & ~n_26486;
assign n_26488 = ~n_26485 & ~n_26487;
assign n_26489 = ~n_26332 & ~n_26488;
assign n_26490 =  n_26332 &  n_26488;
assign n_26491 = ~x_1234 & ~n_26490;
assign n_26492 = ~n_26489 & ~n_26491;
assign n_26493 = ~n_26328 & ~n_26492;
assign n_26494 =  n_26328 &  n_26492;
assign n_26495 = ~x_1233 & ~n_26494;
assign n_26496 = ~n_26493 & ~n_26495;
assign n_26497 = ~n_26326 & ~n_26496;
assign n_26498 =  n_26326 &  n_26496;
assign n_26499 = ~x_1232 & ~n_26498;
assign n_26500 = ~n_26497 & ~n_26499;
assign n_26501 = ~n_26322 & ~n_26500;
assign n_26502 =  n_26322 &  n_26500;
assign n_26503 = ~x_1231 & ~n_26502;
assign n_26504 = ~n_26501 & ~n_26503;
assign n_26505 = ~n_26320 & ~n_26504;
assign n_26506 =  n_26320 &  n_26504;
assign n_26507 = ~x_1230 & ~n_26506;
assign n_26508 = ~n_26505 & ~n_26507;
assign n_26509 = ~n_26316 & ~n_26508;
assign n_26510 =  n_26316 &  n_26508;
assign n_26511 = ~x_1229 & ~n_26510;
assign n_26512 = ~n_26509 & ~n_26511;
assign n_26513 = ~n_26314 & ~n_26512;
assign n_26514 =  n_26314 &  n_26512;
assign n_26515 = ~n_26513 & ~n_26514;
assign n_26516 = ~x_1228 & ~n_26515;
assign n_26517 =  x_1228 &  n_26515;
assign n_26518 = ~n_26516 & ~n_26517;
assign n_26519 = ~n_26509 & ~n_26510;
assign n_26520 =  x_1229 &  n_26519;
assign n_26521 = ~x_1229 & ~n_26519;
assign n_26522 = ~n_26520 & ~n_26521;
assign n_26523 = ~n_26505 & ~n_26506;
assign n_26524 =  x_1230 &  n_26523;
assign n_26525 = ~x_1230 & ~n_26523;
assign n_26526 = ~n_26524 & ~n_26525;
assign n_26527 = ~n_26501 & ~n_26502;
assign n_26528 =  x_1231 &  n_26527;
assign n_26529 = ~x_1231 & ~n_26527;
assign n_26530 = ~n_26528 & ~n_26529;
assign n_26531 = ~n_26497 & ~n_26498;
assign n_26532 =  x_1232 &  n_26531;
assign n_26533 = ~x_1232 & ~n_26531;
assign n_26534 = ~n_26532 & ~n_26533;
assign n_26535 = ~n_26493 & ~n_26494;
assign n_26536 =  x_1233 &  n_26535;
assign n_26537 = ~x_1233 & ~n_26535;
assign n_26538 = ~n_26536 & ~n_26537;
assign n_26539 = ~n_26489 & ~n_26490;
assign n_26540 =  x_1234 &  n_26539;
assign n_26541 = ~x_1234 & ~n_26539;
assign n_26542 = ~n_26540 & ~n_26541;
assign n_26543 = ~n_26485 & ~n_26486;
assign n_26544 =  x_1235 &  n_26543;
assign n_26545 = ~x_1235 & ~n_26543;
assign n_26546 = ~n_26544 & ~n_26545;
assign n_26547 = ~n_26481 & ~n_26482;
assign n_26548 =  x_1236 &  n_26547;
assign n_26549 = ~x_1236 & ~n_26547;
assign n_26550 = ~n_26548 & ~n_26549;
assign n_26551 = ~n_26477 & ~n_26478;
assign n_26552 =  x_1237 &  n_26551;
assign n_26553 = ~x_1237 & ~n_26551;
assign n_26554 = ~n_26552 & ~n_26553;
assign n_26555 = ~n_26473 & ~n_26474;
assign n_26556 =  x_1238 &  n_26555;
assign n_26557 = ~x_1238 & ~n_26555;
assign n_26558 = ~n_26556 & ~n_26557;
assign n_26559 = ~n_26469 & ~n_26470;
assign n_26560 =  x_1239 &  n_26559;
assign n_26561 = ~x_1239 & ~n_26559;
assign n_26562 = ~n_26560 & ~n_26561;
assign n_26563 = ~n_26465 & ~n_26466;
assign n_26564 =  x_1240 &  n_26563;
assign n_26565 = ~x_1240 & ~n_26563;
assign n_26566 = ~n_26564 & ~n_26565;
assign n_26567 = ~n_26461 & ~n_26462;
assign n_26568 =  x_1241 &  n_26567;
assign n_26569 = ~x_1241 & ~n_26567;
assign n_26570 = ~n_26568 & ~n_26569;
assign n_26571 = ~n_26457 & ~n_26458;
assign n_26572 =  x_1242 &  n_26571;
assign n_26573 = ~x_1242 & ~n_26571;
assign n_26574 = ~n_26572 & ~n_26573;
assign n_26575 = ~n_26453 & ~n_26454;
assign n_26576 =  x_1243 &  n_26575;
assign n_26577 = ~x_1243 & ~n_26575;
assign n_26578 = ~n_26576 & ~n_26577;
assign n_26579 = ~n_26449 & ~n_26450;
assign n_26580 =  x_1244 &  n_26579;
assign n_26581 = ~x_1244 & ~n_26579;
assign n_26582 = ~n_26580 & ~n_26581;
assign n_26583 = ~n_26445 & ~n_26446;
assign n_26584 =  x_1245 &  n_26583;
assign n_26585 = ~x_1245 & ~n_26583;
assign n_26586 = ~n_26584 & ~n_26585;
assign n_26587 = ~n_26441 & ~n_26442;
assign n_26588 =  x_1246 &  n_26587;
assign n_26589 = ~x_1246 & ~n_26587;
assign n_26590 = ~n_26588 & ~n_26589;
assign n_26591 = ~n_26437 & ~n_26438;
assign n_26592 =  x_1247 &  n_26591;
assign n_26593 = ~x_1247 & ~n_26591;
assign n_26594 = ~n_26592 & ~n_26593;
assign n_26595 = ~n_26433 & ~n_26434;
assign n_26596 =  x_1248 &  n_26595;
assign n_26597 = ~x_1248 & ~n_26595;
assign n_26598 = ~n_26596 & ~n_26597;
assign n_26599 = ~n_26429 & ~n_26430;
assign n_26600 =  x_1249 &  n_26599;
assign n_26601 = ~x_1249 & ~n_26599;
assign n_26602 = ~n_26600 & ~n_26601;
assign n_26603 = ~n_26425 & ~n_26426;
assign n_26604 =  x_1250 &  n_26603;
assign n_26605 = ~x_1250 & ~n_26603;
assign n_26606 = ~n_26604 & ~n_26605;
assign n_26607 = ~n_26421 & ~n_26422;
assign n_26608 =  x_1251 &  n_26607;
assign n_26609 = ~x_1251 & ~n_26607;
assign n_26610 = ~n_26608 & ~n_26609;
assign n_26611 = ~n_26417 & ~n_26418;
assign n_26612 =  x_1252 &  n_26611;
assign n_26613 = ~x_1252 & ~n_26611;
assign n_26614 = ~n_26612 & ~n_26613;
assign n_26615 = ~n_26413 & ~n_26414;
assign n_26616 =  x_1253 &  n_26615;
assign n_26617 = ~x_1253 & ~n_26615;
assign n_26618 = ~n_26616 & ~n_26617;
assign n_26619 = ~n_26409 & ~n_26410;
assign n_26620 =  x_1254 &  n_26619;
assign n_26621 = ~x_1254 & ~n_26619;
assign n_26622 = ~n_26620 & ~n_26621;
assign n_26623 = ~n_26403 & ~n_26404;
assign n_26624 =  x_1255 &  n_26623;
assign n_26625 = ~x_1255 & ~n_26623;
assign n_26626 = ~n_26624 & ~n_26625;
assign n_26627 = ~n_26396 & ~n_26400;
assign n_26628 = ~n_26399 & ~n_26627;
assign n_26629 = ~n_26396 &  n_26401;
assign n_26630 = ~n_26391 & ~n_26393;
assign n_26631 = ~x_1258 &  x_1290;
assign n_26632 = ~n_26392 & ~n_26631;
assign n_26633 = ~n_26630 &  n_26632;
assign n_26634 = ~n_26629 &  n_26633;
assign n_26635 = ~n_26628 &  n_26634;
assign n_26636 = ~n_26626 &  n_26635;
assign n_26637 = ~n_26622 &  n_26636;
assign n_26638 = ~n_26618 &  n_26637;
assign n_26639 = ~n_26614 &  n_26638;
assign n_26640 = ~n_26610 &  n_26639;
assign n_26641 = ~n_26606 &  n_26640;
assign n_26642 = ~n_26602 &  n_26641;
assign n_26643 = ~n_26598 &  n_26642;
assign n_26644 = ~n_26594 &  n_26643;
assign n_26645 = ~n_26590 &  n_26644;
assign n_26646 = ~n_26586 &  n_26645;
assign n_26647 = ~n_26582 &  n_26646;
assign n_26648 = ~n_26578 &  n_26647;
assign n_26649 = ~n_26574 &  n_26648;
assign n_26650 = ~n_26570 &  n_26649;
assign n_26651 = ~n_26566 &  n_26650;
assign n_26652 = ~n_26562 &  n_26651;
assign n_26653 = ~n_26558 &  n_26652;
assign n_26654 = ~n_26554 &  n_26653;
assign n_26655 = ~n_26550 &  n_26654;
assign n_26656 = ~n_26546 &  n_26655;
assign n_26657 = ~n_26542 &  n_26656;
assign n_26658 = ~n_26538 &  n_26657;
assign n_26659 = ~n_26534 &  n_26658;
assign n_26660 = ~n_26530 &  n_26659;
assign n_26661 = ~n_26526 &  n_26660;
assign n_26662 = ~n_26522 &  n_26661;
assign n_26663 = ~n_26518 &  n_26662;
assign n_26664 = ~x_1259 & ~n_26310;
assign n_26665 =  x_1259 &  n_26310;
assign n_26666 = ~n_26664 & ~n_26665;
assign n_26667 = ~n_26309 &  n_26666;
assign n_26668 =  n_26309 & ~n_26666;
assign n_26669 = ~n_26667 & ~n_26668;
assign n_26670 = ~x_1228 & ~n_26514;
assign n_26671 = ~n_26513 & ~n_26670;
assign n_26672 =  n_26669 &  n_26671;
assign n_26673 = ~n_26669 & ~n_26671;
assign n_26674 = ~n_26672 & ~n_26673;
assign n_26675 =  x_1227 & ~n_26674;
assign n_26676 = ~x_1227 &  n_26674;
assign n_26677 = ~n_26675 & ~n_26676;
assign n_26678 =  n_26663 &  n_26677;
assign n_26679 =  n_26229 &  n_26678;
assign n_26680 = ~x_2280 & ~x_2281;
assign n_26681 = ~x_2279 &  n_26680;
assign n_26682 = ~x_2278 &  n_26681;
assign n_26683 = ~x_2277 & ~x_2282;
assign n_26684 =  n_26682 &  n_26683;
assign n_26685 = ~x_2276 &  n_26684;
assign n_26686 = ~x_2275 &  n_26685;
assign n_26687 = ~x_2274 &  n_26686;
assign n_26688 = ~x_2273 &  n_26687;
assign n_26689 = ~x_2272 &  n_26688;
assign n_26690 = ~x_2271 &  n_26689;
assign n_26691 = ~x_2270 &  n_26690;
assign n_26692 = ~x_2269 &  n_26691;
assign n_26693 = ~x_2268 &  n_26692;
assign n_26694 = ~x_2267 &  n_26693;
assign n_26695 = ~x_2266 &  n_26694;
assign n_26696 = ~x_2265 &  n_26695;
assign n_26697 = ~x_2264 &  n_26696;
assign n_26698 = ~x_2263 &  n_26697;
assign n_26699 = ~x_2262 &  n_26698;
assign n_26700 = ~x_2261 &  n_26699;
assign n_26701 = ~x_2260 &  n_26700;
assign n_26702 = ~x_2259 &  n_26701;
assign n_26703 = ~x_2258 &  n_26702;
assign n_26704 = ~x_2257 &  n_26703;
assign n_26705 = ~x_2256 &  n_26704;
assign n_26706 = ~x_2255 &  n_26705;
assign n_26707 = ~x_2254 &  n_26706;
assign n_26708 = ~x_2253 &  n_26707;
assign n_26709 =  x_2253 & ~n_26707;
assign n_26710 = ~n_26708 & ~n_26709;
assign n_26711 =  x_2255 & ~n_26705;
assign n_26712 = ~n_26706 & ~n_26711;
assign n_26713 =  x_2257 & ~n_26703;
assign n_26714 = ~n_26704 & ~n_26713;
assign n_26715 =  x_2259 & ~n_26701;
assign n_26716 = ~n_26702 & ~n_26715;
assign n_26717 =  x_2261 & ~n_26699;
assign n_26718 = ~n_26700 & ~n_26717;
assign n_26719 =  x_2263 & ~n_26697;
assign n_26720 = ~n_26698 & ~n_26719;
assign n_26721 =  x_2265 & ~n_26695;
assign n_26722 = ~n_26696 & ~n_26721;
assign n_26723 =  x_2267 & ~n_26693;
assign n_26724 = ~n_26694 & ~n_26723;
assign n_26725 =  x_2269 & ~n_26691;
assign n_26726 = ~n_26692 & ~n_26725;
assign n_26727 =  x_2271 & ~n_26689;
assign n_26728 = ~n_26690 & ~n_26727;
assign n_26729 =  x_2273 & ~n_26687;
assign n_26730 = ~n_26688 & ~n_26729;
assign n_26731 =  x_2275 & ~n_26685;
assign n_26732 = ~n_26686 & ~n_26731;
assign n_26733 = ~x_2277 &  x_2282;
assign n_26734 =  n_26682 &  n_26733;
assign n_26735 = ~x_2276 &  n_26734;
assign n_26736 =  n_26732 &  n_26735;
assign n_26737 = ~x_2274 &  n_26736;
assign n_26738 =  n_26730 &  n_26737;
assign n_26739 = ~x_2272 &  n_26738;
assign n_26740 =  n_26728 &  n_26739;
assign n_26741 = ~x_2270 &  n_26740;
assign n_26742 =  n_26726 &  n_26741;
assign n_26743 = ~x_2268 &  n_26742;
assign n_26744 =  n_26724 &  n_26743;
assign n_26745 = ~x_2266 &  n_26744;
assign n_26746 =  n_26722 &  n_26745;
assign n_26747 = ~x_2264 &  n_26746;
assign n_26748 =  n_26720 &  n_26747;
assign n_26749 = ~x_2262 &  n_26748;
assign n_26750 =  n_26718 &  n_26749;
assign n_26751 = ~x_2260 &  n_26750;
assign n_26752 =  n_26716 &  n_26751;
assign n_26753 = ~x_2258 &  n_26752;
assign n_26754 =  n_26714 &  n_26753;
assign n_26755 = ~x_2256 &  n_26754;
assign n_26756 =  n_26712 &  n_26755;
assign n_26757 = ~x_2254 &  n_26756;
assign n_26758 =  n_26710 &  n_26757;
assign n_26759 = ~x_2252 &  n_26758;
assign n_26760 = ~x_2252 &  n_26708;
assign n_26761 = ~x_2251 & ~n_26760;
assign n_26762 =  x_2251 &  n_26760;
assign n_26763 = ~n_26761 & ~n_26762;
assign n_26764 = ~n_26759 &  n_26763;
assign n_26765 =  n_26759 & ~n_26763;
assign n_26766 = ~n_26764 & ~n_26765;
assign n_26767 =  x_2252 & ~n_26708;
assign n_26768 = ~n_26760 & ~n_26767;
assign n_26769 = ~n_26758 & ~n_26768;
assign n_26770 = ~n_26759 & ~n_26769;
assign n_26771 = ~n_26710 & ~n_26757;
assign n_26772 = ~n_26758 & ~n_26771;
assign n_26773 =  x_2254 & ~n_26706;
assign n_26774 = ~n_26707 & ~n_26773;
assign n_26775 = ~n_26756 & ~n_26774;
assign n_26776 = ~n_26757 & ~n_26775;
assign n_26777 = ~n_26712 & ~n_26755;
assign n_26778 = ~n_26756 & ~n_26777;
assign n_26779 =  x_2256 & ~n_26704;
assign n_26780 = ~n_26705 & ~n_26779;
assign n_26781 = ~n_26754 & ~n_26780;
assign n_26782 = ~n_26755 & ~n_26781;
assign n_26783 = ~n_26714 & ~n_26753;
assign n_26784 = ~n_26754 & ~n_26783;
assign n_26785 =  x_2258 & ~n_26702;
assign n_26786 = ~n_26703 & ~n_26785;
assign n_26787 = ~n_26752 & ~n_26786;
assign n_26788 = ~n_26753 & ~n_26787;
assign n_26789 = ~n_26716 & ~n_26751;
assign n_26790 = ~n_26752 & ~n_26789;
assign n_26791 =  x_2260 & ~n_26700;
assign n_26792 = ~n_26701 & ~n_26791;
assign n_26793 = ~n_26750 & ~n_26792;
assign n_26794 = ~n_26751 & ~n_26793;
assign n_26795 = ~n_26718 & ~n_26749;
assign n_26796 = ~n_26750 & ~n_26795;
assign n_26797 =  x_2262 & ~n_26698;
assign n_26798 = ~n_26699 & ~n_26797;
assign n_26799 = ~n_26748 & ~n_26798;
assign n_26800 = ~n_26749 & ~n_26799;
assign n_26801 = ~n_26720 & ~n_26747;
assign n_26802 = ~n_26748 & ~n_26801;
assign n_26803 =  x_2264 & ~n_26696;
assign n_26804 = ~n_26697 & ~n_26803;
assign n_26805 = ~n_26746 & ~n_26804;
assign n_26806 = ~n_26747 & ~n_26805;
assign n_26807 = ~n_26722 & ~n_26745;
assign n_26808 = ~n_26746 & ~n_26807;
assign n_26809 =  x_2266 & ~n_26694;
assign n_26810 = ~n_26695 & ~n_26809;
assign n_26811 = ~n_26744 & ~n_26810;
assign n_26812 = ~n_26745 & ~n_26811;
assign n_26813 = ~n_26724 & ~n_26743;
assign n_26814 = ~n_26744 & ~n_26813;
assign n_26815 =  x_2268 & ~n_26692;
assign n_26816 = ~n_26693 & ~n_26815;
assign n_26817 = ~n_26742 & ~n_26816;
assign n_26818 = ~n_26743 & ~n_26817;
assign n_26819 = ~n_26726 & ~n_26741;
assign n_26820 = ~n_26742 & ~n_26819;
assign n_26821 =  x_2270 & ~n_26690;
assign n_26822 = ~n_26691 & ~n_26821;
assign n_26823 = ~n_26740 & ~n_26822;
assign n_26824 = ~n_26741 & ~n_26823;
assign n_26825 = ~n_26728 & ~n_26739;
assign n_26826 = ~n_26740 & ~n_26825;
assign n_26827 =  x_2272 & ~n_26688;
assign n_26828 = ~n_26689 & ~n_26827;
assign n_26829 = ~n_26738 & ~n_26828;
assign n_26830 = ~n_26739 & ~n_26829;
assign n_26831 = ~n_26730 & ~n_26737;
assign n_26832 = ~n_26738 & ~n_26831;
assign n_26833 =  x_2274 & ~n_26686;
assign n_26834 = ~n_26687 & ~n_26833;
assign n_26835 = ~n_26736 & ~n_26834;
assign n_26836 = ~n_26737 & ~n_26835;
assign n_26837 = ~n_26732 & ~n_26735;
assign n_26838 = ~n_26736 & ~n_26837;
assign n_26839 = ~n_26684 & ~n_26734;
assign n_26840 =  x_2276 & ~n_26839;
assign n_26841 = ~x_2276 &  n_26839;
assign n_26842 = ~n_26840 & ~n_26841;
assign n_26843 =  x_2277 & ~n_26682;
assign n_26844 =  n_26839 & ~n_26843;
assign n_26845 =  x_2279 & ~n_26680;
assign n_26846 = ~n_26681 & ~n_26845;
assign n_26847 = ~x_1801 & ~x_2281;
assign n_26848 =  x_1802 & ~x_2282;
assign n_26849 =  x_1801 &  x_2281;
assign n_26850 = ~n_26848 & ~n_26849;
assign n_26851 = ~n_26847 & ~n_26850;
assign n_26852 =  x_2280 &  x_2281;
assign n_26853 = ~n_26680 & ~n_26852;
assign n_26854 =  x_1800 &  n_26853;
assign n_26855 = ~n_26851 & ~n_26854;
assign n_26856 = ~x_1800 & ~n_26853;
assign n_26857 = ~n_26855 & ~n_26856;
assign n_26858 = ~n_26846 & ~n_26857;
assign n_26859 =  n_26846 &  n_26857;
assign n_26860 = ~x_1799 & ~n_26859;
assign n_26861 = ~n_26858 & ~n_26860;
assign n_26862 =  x_2278 & ~n_26681;
assign n_26863 = ~n_26682 & ~n_26862;
assign n_26864 = ~n_26861 & ~n_26863;
assign n_26865 =  n_26861 &  n_26863;
assign n_26866 = ~x_1798 & ~n_26865;
assign n_26867 = ~n_26864 & ~n_26866;
assign n_26868 = ~n_26844 & ~n_26867;
assign n_26869 =  n_26844 &  n_26867;
assign n_26870 = ~x_1797 & ~n_26869;
assign n_26871 = ~n_26868 & ~n_26870;
assign n_26872 =  n_26842 & ~n_26871;
assign n_26873 = ~n_26842 &  n_26871;
assign n_26874 = ~x_1796 & ~n_26873;
assign n_26875 = ~n_26872 & ~n_26874;
assign n_26876 = ~n_26838 & ~n_26875;
assign n_26877 =  n_26838 &  n_26875;
assign n_26878 = ~x_1795 & ~n_26877;
assign n_26879 = ~n_26876 & ~n_26878;
assign n_26880 = ~n_26836 & ~n_26879;
assign n_26881 =  n_26836 &  n_26879;
assign n_26882 = ~x_1794 & ~n_26881;
assign n_26883 = ~n_26880 & ~n_26882;
assign n_26884 = ~n_26832 & ~n_26883;
assign n_26885 =  n_26832 &  n_26883;
assign n_26886 = ~x_1793 & ~n_26885;
assign n_26887 = ~n_26884 & ~n_26886;
assign n_26888 = ~n_26830 & ~n_26887;
assign n_26889 =  n_26830 &  n_26887;
assign n_26890 = ~x_1792 & ~n_26889;
assign n_26891 = ~n_26888 & ~n_26890;
assign n_26892 = ~n_26826 & ~n_26891;
assign n_26893 =  n_26826 &  n_26891;
assign n_26894 = ~x_1791 & ~n_26893;
assign n_26895 = ~n_26892 & ~n_26894;
assign n_26896 = ~n_26824 & ~n_26895;
assign n_26897 =  n_26824 &  n_26895;
assign n_26898 = ~x_1790 & ~n_26897;
assign n_26899 = ~n_26896 & ~n_26898;
assign n_26900 = ~n_26820 & ~n_26899;
assign n_26901 =  n_26820 &  n_26899;
assign n_26902 = ~x_1789 & ~n_26901;
assign n_26903 = ~n_26900 & ~n_26902;
assign n_26904 = ~n_26818 & ~n_26903;
assign n_26905 =  n_26818 &  n_26903;
assign n_26906 = ~x_1788 & ~n_26905;
assign n_26907 = ~n_26904 & ~n_26906;
assign n_26908 = ~n_26814 & ~n_26907;
assign n_26909 =  n_26814 &  n_26907;
assign n_26910 = ~x_1787 & ~n_26909;
assign n_26911 = ~n_26908 & ~n_26910;
assign n_26912 = ~n_26812 & ~n_26911;
assign n_26913 =  n_26812 &  n_26911;
assign n_26914 = ~x_1786 & ~n_26913;
assign n_26915 = ~n_26912 & ~n_26914;
assign n_26916 = ~n_26808 & ~n_26915;
assign n_26917 =  n_26808 &  n_26915;
assign n_26918 = ~x_1785 & ~n_26917;
assign n_26919 = ~n_26916 & ~n_26918;
assign n_26920 = ~n_26806 & ~n_26919;
assign n_26921 =  n_26806 &  n_26919;
assign n_26922 = ~x_1784 & ~n_26921;
assign n_26923 = ~n_26920 & ~n_26922;
assign n_26924 = ~n_26802 & ~n_26923;
assign n_26925 =  n_26802 &  n_26923;
assign n_26926 = ~x_1783 & ~n_26925;
assign n_26927 = ~n_26924 & ~n_26926;
assign n_26928 = ~n_26800 & ~n_26927;
assign n_26929 =  n_26800 &  n_26927;
assign n_26930 = ~x_1782 & ~n_26929;
assign n_26931 = ~n_26928 & ~n_26930;
assign n_26932 = ~n_26796 & ~n_26931;
assign n_26933 =  n_26796 &  n_26931;
assign n_26934 = ~x_1781 & ~n_26933;
assign n_26935 = ~n_26932 & ~n_26934;
assign n_26936 = ~n_26794 & ~n_26935;
assign n_26937 =  n_26794 &  n_26935;
assign n_26938 = ~x_1780 & ~n_26937;
assign n_26939 = ~n_26936 & ~n_26938;
assign n_26940 = ~n_26790 & ~n_26939;
assign n_26941 =  n_26790 &  n_26939;
assign n_26942 = ~x_1779 & ~n_26941;
assign n_26943 = ~n_26940 & ~n_26942;
assign n_26944 = ~n_26788 & ~n_26943;
assign n_26945 =  n_26788 &  n_26943;
assign n_26946 = ~x_1778 & ~n_26945;
assign n_26947 = ~n_26944 & ~n_26946;
assign n_26948 = ~n_26784 & ~n_26947;
assign n_26949 =  n_26784 &  n_26947;
assign n_26950 = ~x_1777 & ~n_26949;
assign n_26951 = ~n_26948 & ~n_26950;
assign n_26952 = ~n_26782 & ~n_26951;
assign n_26953 =  n_26782 &  n_26951;
assign n_26954 = ~x_1776 & ~n_26953;
assign n_26955 = ~n_26952 & ~n_26954;
assign n_26956 = ~n_26778 & ~n_26955;
assign n_26957 =  n_26778 &  n_26955;
assign n_26958 = ~x_1775 & ~n_26957;
assign n_26959 = ~n_26956 & ~n_26958;
assign n_26960 = ~n_26776 & ~n_26959;
assign n_26961 =  n_26776 &  n_26959;
assign n_26962 = ~x_1774 & ~n_26961;
assign n_26963 = ~n_26960 & ~n_26962;
assign n_26964 = ~n_26772 & ~n_26963;
assign n_26965 =  n_26772 &  n_26963;
assign n_26966 = ~x_1773 & ~n_26965;
assign n_26967 = ~n_26964 & ~n_26966;
assign n_26968 = ~n_26770 & ~n_26967;
assign n_26969 =  n_26770 &  n_26967;
assign n_26970 = ~x_1772 & ~n_26969;
assign n_26971 = ~n_26968 & ~n_26970;
assign n_26972 =  n_26766 &  n_26971;
assign n_26973 = ~n_26766 & ~n_26971;
assign n_26974 = ~n_26972 & ~n_26973;
assign n_26975 = ~x_1771 & ~n_26974;
assign n_26976 =  x_1771 &  n_26974;
assign n_26977 = ~n_26975 & ~n_26976;
assign n_26978 = ~n_26968 & ~n_26969;
assign n_26979 =  x_1772 &  n_26978;
assign n_26980 = ~x_1772 & ~n_26978;
assign n_26981 = ~n_26979 & ~n_26980;
assign n_26982 = ~n_26964 & ~n_26965;
assign n_26983 =  x_1773 &  n_26982;
assign n_26984 = ~x_1773 & ~n_26982;
assign n_26985 = ~n_26983 & ~n_26984;
assign n_26986 = ~n_26960 & ~n_26961;
assign n_26987 =  x_1774 &  n_26986;
assign n_26988 = ~x_1774 & ~n_26986;
assign n_26989 = ~n_26987 & ~n_26988;
assign n_26990 = ~n_26956 & ~n_26957;
assign n_26991 =  x_1775 &  n_26990;
assign n_26992 = ~x_1775 & ~n_26990;
assign n_26993 = ~n_26991 & ~n_26992;
assign n_26994 = ~n_26952 & ~n_26953;
assign n_26995 =  x_1776 &  n_26994;
assign n_26996 = ~x_1776 & ~n_26994;
assign n_26997 = ~n_26995 & ~n_26996;
assign n_26998 = ~n_26948 & ~n_26949;
assign n_26999 =  x_1777 &  n_26998;
assign n_27000 = ~x_1777 & ~n_26998;
assign n_27001 = ~n_26999 & ~n_27000;
assign n_27002 = ~n_26944 & ~n_26945;
assign n_27003 =  x_1778 &  n_27002;
assign n_27004 = ~x_1778 & ~n_27002;
assign n_27005 = ~n_27003 & ~n_27004;
assign n_27006 = ~n_26940 & ~n_26941;
assign n_27007 =  x_1779 &  n_27006;
assign n_27008 = ~x_1779 & ~n_27006;
assign n_27009 = ~n_27007 & ~n_27008;
assign n_27010 = ~n_26936 & ~n_26937;
assign n_27011 =  x_1780 &  n_27010;
assign n_27012 = ~x_1780 & ~n_27010;
assign n_27013 = ~n_27011 & ~n_27012;
assign n_27014 = ~n_26932 & ~n_26933;
assign n_27015 =  x_1781 &  n_27014;
assign n_27016 = ~x_1781 & ~n_27014;
assign n_27017 = ~n_27015 & ~n_27016;
assign n_27018 = ~n_26928 & ~n_26929;
assign n_27019 =  x_1782 &  n_27018;
assign n_27020 = ~x_1782 & ~n_27018;
assign n_27021 = ~n_27019 & ~n_27020;
assign n_27022 = ~n_26924 & ~n_26925;
assign n_27023 =  x_1783 &  n_27022;
assign n_27024 = ~x_1783 & ~n_27022;
assign n_27025 = ~n_27023 & ~n_27024;
assign n_27026 = ~n_26920 & ~n_26921;
assign n_27027 =  x_1784 &  n_27026;
assign n_27028 = ~x_1784 & ~n_27026;
assign n_27029 = ~n_27027 & ~n_27028;
assign n_27030 = ~n_26916 & ~n_26917;
assign n_27031 =  x_1785 &  n_27030;
assign n_27032 = ~x_1785 & ~n_27030;
assign n_27033 = ~n_27031 & ~n_27032;
assign n_27034 = ~n_26912 & ~n_26913;
assign n_27035 =  x_1786 &  n_27034;
assign n_27036 = ~x_1786 & ~n_27034;
assign n_27037 = ~n_27035 & ~n_27036;
assign n_27038 = ~n_26908 & ~n_26909;
assign n_27039 =  x_1787 &  n_27038;
assign n_27040 = ~x_1787 & ~n_27038;
assign n_27041 = ~n_27039 & ~n_27040;
assign n_27042 = ~n_26904 & ~n_26905;
assign n_27043 =  x_1788 &  n_27042;
assign n_27044 = ~x_1788 & ~n_27042;
assign n_27045 = ~n_27043 & ~n_27044;
assign n_27046 = ~n_26900 & ~n_26901;
assign n_27047 =  x_1789 &  n_27046;
assign n_27048 = ~x_1789 & ~n_27046;
assign n_27049 = ~n_27047 & ~n_27048;
assign n_27050 = ~n_26896 & ~n_26897;
assign n_27051 =  x_1790 &  n_27050;
assign n_27052 = ~x_1790 & ~n_27050;
assign n_27053 = ~n_27051 & ~n_27052;
assign n_27054 = ~n_26892 & ~n_26893;
assign n_27055 =  x_1791 &  n_27054;
assign n_27056 = ~x_1791 & ~n_27054;
assign n_27057 = ~n_27055 & ~n_27056;
assign n_27058 = ~n_26888 & ~n_26889;
assign n_27059 =  x_1792 &  n_27058;
assign n_27060 = ~x_1792 & ~n_27058;
assign n_27061 = ~n_27059 & ~n_27060;
assign n_27062 = ~n_26884 & ~n_26885;
assign n_27063 =  x_1793 &  n_27062;
assign n_27064 = ~x_1793 & ~n_27062;
assign n_27065 = ~n_27063 & ~n_27064;
assign n_27066 = ~n_26880 & ~n_26881;
assign n_27067 =  x_1794 &  n_27066;
assign n_27068 = ~x_1794 & ~n_27066;
assign n_27069 = ~n_27067 & ~n_27068;
assign n_27070 = ~n_26876 & ~n_26877;
assign n_27071 =  x_1795 &  n_27070;
assign n_27072 = ~x_1795 & ~n_27070;
assign n_27073 = ~n_27071 & ~n_27072;
assign n_27074 = ~n_26872 & ~n_26873;
assign n_27075 =  x_1796 &  n_27074;
assign n_27076 = ~x_1796 & ~n_27074;
assign n_27077 = ~n_27075 & ~n_27076;
assign n_27078 = ~n_26868 & ~n_26869;
assign n_27079 =  x_1797 &  n_27078;
assign n_27080 = ~x_1797 & ~n_27078;
assign n_27081 = ~n_27079 & ~n_27080;
assign n_27082 = ~n_26864 & ~n_26865;
assign n_27083 =  x_1798 &  n_27082;
assign n_27084 = ~x_1798 & ~n_27082;
assign n_27085 = ~n_27083 & ~n_27084;
assign n_27086 = ~n_26858 & ~n_26859;
assign n_27087 =  x_1799 &  n_27086;
assign n_27088 = ~x_1799 & ~n_27086;
assign n_27089 = ~n_27087 & ~n_27088;
assign n_27090 = ~n_26847 & ~n_26849;
assign n_27091 =  x_1800 &  x_2280;
assign n_27092 = ~x_1800 & ~x_2280;
assign n_27093 = ~n_27091 & ~n_27092;
assign n_27094 =  x_1802 &  x_2282;
assign n_27095 = ~x_1802 & ~x_2282;
assign n_27096 = ~n_27094 & ~n_27095;
assign n_27097 = ~n_27093 & ~n_27096;
assign n_27098 = ~n_27090 &  n_27097;
assign n_27099 =  n_8060 &  n_27098;
assign n_27100 =  n_588 &  n_27099;
assign n_27101 = ~n_27089 &  n_27100;
assign n_27102 = ~n_27085 &  n_27101;
assign n_27103 = ~n_27081 &  n_27102;
assign n_27104 = ~n_27077 &  n_27103;
assign n_27105 = ~n_27073 &  n_27104;
assign n_27106 = ~n_27069 &  n_27105;
assign n_27107 = ~n_27065 &  n_27106;
assign n_27108 = ~n_27061 &  n_27107;
assign n_27109 = ~n_27057 &  n_27108;
assign n_27110 = ~n_27053 &  n_27109;
assign n_27111 = ~n_27049 &  n_27110;
assign n_27112 = ~n_27045 &  n_27111;
assign n_27113 = ~n_27041 &  n_27112;
assign n_27114 = ~n_27037 &  n_27113;
assign n_27115 = ~n_27033 &  n_27114;
assign n_27116 = ~n_27029 &  n_27115;
assign n_27117 = ~n_27025 &  n_27116;
assign n_27118 = ~n_27021 &  n_27117;
assign n_27119 = ~n_27017 &  n_27118;
assign n_27120 = ~n_27013 &  n_27119;
assign n_27121 = ~n_27009 &  n_27120;
assign n_27122 = ~n_27005 &  n_27121;
assign n_27123 = ~n_27001 &  n_27122;
assign n_27124 = ~n_26997 &  n_27123;
assign n_27125 = ~n_26993 &  n_27124;
assign n_27126 = ~n_26989 &  n_27125;
assign n_27127 = ~n_26985 &  n_27126;
assign n_27128 = ~n_26981 &  n_27127;
assign n_27129 = ~n_26977 &  n_27128;
assign n_27130 = ~x_1547 &  x_2187;
assign n_27131 =  x_1547 & ~x_2187;
assign n_27132 =  x_1548 & ~x_2188;
assign n_27133 = ~x_1548 &  x_2188;
assign n_27134 =  x_1549 & ~x_2189;
assign n_27135 = ~x_1549 &  x_2189;
assign n_27136 =  x_1550 & ~x_2190;
assign n_27137 = ~x_1550 &  x_2190;
assign n_27138 =  x_1551 & ~x_2191;
assign n_27139 = ~x_1551 &  x_2191;
assign n_27140 =  x_1552 & ~x_2192;
assign n_27141 = ~x_1552 &  x_2192;
assign n_27142 =  x_1553 & ~x_2193;
assign n_27143 = ~x_1553 &  x_2193;
assign n_27144 =  x_1554 & ~x_2194;
assign n_27145 = ~x_1554 &  x_2194;
assign n_27146 =  x_1555 & ~x_2195;
assign n_27147 = ~x_1555 &  x_2195;
assign n_27148 =  x_1556 & ~x_2196;
assign n_27149 = ~x_1556 &  x_2196;
assign n_27150 =  x_1557 & ~x_2197;
assign n_27151 = ~x_1557 &  x_2197;
assign n_27152 =  x_1558 & ~x_2198;
assign n_27153 = ~x_1558 &  x_2198;
assign n_27154 =  x_1559 & ~x_2199;
assign n_27155 = ~x_1559 &  x_2199;
assign n_27156 =  x_1560 & ~x_2200;
assign n_27157 = ~x_1560 &  x_2200;
assign n_27158 =  x_1561 & ~x_2201;
assign n_27159 = ~x_1561 &  x_2201;
assign n_27160 =  x_1562 & ~x_2202;
assign n_27161 = ~x_1562 &  x_2202;
assign n_27162 =  x_1563 & ~x_2203;
assign n_27163 = ~x_1563 &  x_2203;
assign n_27164 =  x_1564 & ~x_2204;
assign n_27165 = ~x_1564 &  x_2204;
assign n_27166 =  x_1565 & ~x_2205;
assign n_27167 = ~x_1565 &  x_2205;
assign n_27168 =  x_1566 & ~x_2206;
assign n_27169 = ~x_1566 &  x_2206;
assign n_27170 =  x_1567 & ~x_2207;
assign n_27171 = ~x_1567 &  x_2207;
assign n_27172 =  x_1568 & ~x_2208;
assign n_27173 = ~x_1568 &  x_2208;
assign n_27174 =  x_1569 & ~x_2209;
assign n_27175 = ~x_1569 &  x_2209;
assign n_27176 =  x_1570 & ~x_2210;
assign n_27177 = ~x_1570 &  x_2210;
assign n_27178 =  x_1571 & ~x_2211;
assign n_27179 = ~x_1571 &  x_2211;
assign n_27180 =  x_1572 & ~x_2212;
assign n_27181 = ~x_1572 &  x_2212;
assign n_27182 =  x_1573 & ~x_2213;
assign n_27183 = ~x_1573 &  x_2213;
assign n_27184 =  x_1574 & ~x_2214;
assign n_27185 = ~x_1574 &  x_2214;
assign n_27186 =  x_1575 & ~x_2215;
assign n_27187 = ~x_1575 &  x_2215;
assign n_27188 =  x_1577 & ~x_2217;
assign n_27189 = ~x_1577 &  x_2217;
assign n_27190 =  x_1578 & ~x_2218;
assign n_27191 = ~n_27189 &  n_27190;
assign n_27192 = ~n_27188 & ~n_27191;
assign n_27193 =  x_2216 &  n_27192;
assign n_27194 =  x_1576 & ~n_27193;
assign n_27195 = ~x_2216 & ~n_27192;
assign n_27196 = ~n_27194 & ~n_27195;
assign n_27197 = ~n_27187 & ~n_27196;
assign n_27198 = ~n_27186 & ~n_27197;
assign n_27199 = ~n_27185 & ~n_27198;
assign n_27200 = ~n_27184 & ~n_27199;
assign n_27201 = ~n_27183 & ~n_27200;
assign n_27202 = ~n_27182 & ~n_27201;
assign n_27203 = ~n_27181 & ~n_27202;
assign n_27204 = ~n_27180 & ~n_27203;
assign n_27205 = ~n_27179 & ~n_27204;
assign n_27206 = ~n_27178 & ~n_27205;
assign n_27207 = ~n_27177 & ~n_27206;
assign n_27208 = ~n_27176 & ~n_27207;
assign n_27209 = ~n_27175 & ~n_27208;
assign n_27210 = ~n_27174 & ~n_27209;
assign n_27211 = ~n_27173 & ~n_27210;
assign n_27212 = ~n_27172 & ~n_27211;
assign n_27213 = ~n_27171 & ~n_27212;
assign n_27214 = ~n_27170 & ~n_27213;
assign n_27215 = ~n_27169 & ~n_27214;
assign n_27216 = ~n_27168 & ~n_27215;
assign n_27217 = ~n_27167 & ~n_27216;
assign n_27218 = ~n_27166 & ~n_27217;
assign n_27219 = ~n_27165 & ~n_27218;
assign n_27220 = ~n_27164 & ~n_27219;
assign n_27221 = ~n_27163 & ~n_27220;
assign n_27222 = ~n_27162 & ~n_27221;
assign n_27223 = ~n_27161 & ~n_27222;
assign n_27224 = ~n_27160 & ~n_27223;
assign n_27225 = ~n_27159 & ~n_27224;
assign n_27226 = ~n_27158 & ~n_27225;
assign n_27227 = ~n_27157 & ~n_27226;
assign n_27228 = ~n_27156 & ~n_27227;
assign n_27229 = ~n_27155 & ~n_27228;
assign n_27230 = ~n_27154 & ~n_27229;
assign n_27231 = ~n_27153 & ~n_27230;
assign n_27232 = ~n_27152 & ~n_27231;
assign n_27233 = ~n_27151 & ~n_27232;
assign n_27234 = ~n_27150 & ~n_27233;
assign n_27235 = ~n_27149 & ~n_27234;
assign n_27236 = ~n_27148 & ~n_27235;
assign n_27237 = ~n_27147 & ~n_27236;
assign n_27238 = ~n_27146 & ~n_27237;
assign n_27239 = ~n_27145 & ~n_27238;
assign n_27240 = ~n_27144 & ~n_27239;
assign n_27241 = ~n_27143 & ~n_27240;
assign n_27242 = ~n_27142 & ~n_27241;
assign n_27243 = ~n_27141 & ~n_27242;
assign n_27244 = ~n_27140 & ~n_27243;
assign n_27245 = ~n_27139 & ~n_27244;
assign n_27246 = ~n_27138 & ~n_27245;
assign n_27247 = ~n_27137 & ~n_27246;
assign n_27248 = ~n_27136 & ~n_27247;
assign n_27249 = ~n_27135 & ~n_27248;
assign n_27250 = ~n_27134 & ~n_27249;
assign n_27251 = ~n_27133 & ~n_27250;
assign n_27252 = ~n_27132 & ~n_27251;
assign n_27253 = ~n_27131 & ~n_27252;
assign n_27254 = ~n_27130 & ~n_27253;
assign n_27255 =  x_33 & ~x_34;
assign n_27256 = ~x_35 &  n_27255;
assign n_27257 =  x_36 &  n_27256;
assign n_27258 = ~x_37 &  n_27257;
assign n_27259 = ~x_38 &  n_27258;
assign n_27260 =  n_27254 &  n_27259;
assign n_27261 =  n_3664 &  n_27260;
assign n_27262 =  n_27257 &  n_10319;
assign n_27263 =  n_27254 &  n_27262;
assign n_27264 =  n_27263 &  n_10318;
assign n_27265 = ~n_27261 & ~n_27264;
assign n_27266 =  n_27256 &  n_2295;
assign n_27267 = ~x_38 &  n_27266;
assign n_27268 =  n_27254 &  n_27267;
assign n_27269 =  n_3664 &  n_27268;
assign n_27270 =  n_8818 &  n_27268;
assign n_27271 = ~n_27269 & ~n_27270;
assign n_27272 =  n_27265 &  n_27271;
assign n_27273 =  x_36 &  n_6;
assign n_27274 = ~x_37 &  n_27273;
assign n_27275 = ~x_1163 &  x_2187;
assign n_27276 =  x_1163 & ~x_2187;
assign n_27277 =  x_1164 & ~x_2188;
assign n_27278 = ~x_1164 &  x_2188;
assign n_27279 =  x_1165 & ~x_2189;
assign n_27280 = ~x_1165 &  x_2189;
assign n_27281 =  x_1166 & ~x_2190;
assign n_27282 = ~x_1166 &  x_2190;
assign n_27283 =  x_1167 & ~x_2191;
assign n_27284 = ~x_1167 &  x_2191;
assign n_27285 =  x_1168 & ~x_2192;
assign n_27286 = ~x_1168 &  x_2192;
assign n_27287 =  x_1169 & ~x_2193;
assign n_27288 = ~x_1169 &  x_2193;
assign n_27289 =  x_1170 & ~x_2194;
assign n_27290 = ~x_1170 &  x_2194;
assign n_27291 =  x_1171 & ~x_2195;
assign n_27292 = ~x_1171 &  x_2195;
assign n_27293 =  x_1172 & ~x_2196;
assign n_27294 = ~x_1172 &  x_2196;
assign n_27295 =  x_1173 & ~x_2197;
assign n_27296 = ~x_1173 &  x_2197;
assign n_27297 =  x_1174 & ~x_2198;
assign n_27298 = ~x_1174 &  x_2198;
assign n_27299 =  x_1175 & ~x_2199;
assign n_27300 = ~x_1175 &  x_2199;
assign n_27301 =  x_1176 & ~x_2200;
assign n_27302 = ~x_1176 &  x_2200;
assign n_27303 =  x_1177 & ~x_2201;
assign n_27304 = ~x_1177 &  x_2201;
assign n_27305 =  x_1178 & ~x_2202;
assign n_27306 = ~x_1178 &  x_2202;
assign n_27307 =  x_1179 & ~x_2203;
assign n_27308 = ~x_1179 &  x_2203;
assign n_27309 =  x_1180 & ~x_2204;
assign n_27310 = ~x_1180 &  x_2204;
assign n_27311 =  x_1181 & ~x_2205;
assign n_27312 = ~x_1181 &  x_2205;
assign n_27313 =  x_1182 & ~x_2206;
assign n_27314 = ~x_1182 &  x_2206;
assign n_27315 =  x_1183 & ~x_2207;
assign n_27316 = ~x_1183 &  x_2207;
assign n_27317 =  x_1184 & ~x_2208;
assign n_27318 = ~x_1184 &  x_2208;
assign n_27319 =  x_1185 & ~x_2209;
assign n_27320 = ~x_1185 &  x_2209;
assign n_27321 =  x_1186 & ~x_2210;
assign n_27322 = ~x_1186 &  x_2210;
assign n_27323 =  x_1187 & ~x_2211;
assign n_27324 = ~x_1187 &  x_2211;
assign n_27325 =  x_1188 & ~x_2212;
assign n_27326 = ~x_1188 &  x_2212;
assign n_27327 =  x_1189 & ~x_2213;
assign n_27328 = ~x_1189 &  x_2213;
assign n_27329 =  x_1190 & ~x_2214;
assign n_27330 = ~x_1190 &  x_2214;
assign n_27331 =  x_1191 & ~x_2215;
assign n_27332 = ~x_1191 &  x_2215;
assign n_27333 =  x_1193 & ~x_2217;
assign n_27334 = ~x_1193 &  x_2217;
assign n_27335 =  x_1194 & ~x_2218;
assign n_27336 = ~n_27334 &  n_27335;
assign n_27337 = ~n_27333 & ~n_27336;
assign n_27338 =  x_2216 &  n_27337;
assign n_27339 =  x_1192 & ~n_27338;
assign n_27340 = ~x_2216 & ~n_27337;
assign n_27341 = ~n_27339 & ~n_27340;
assign n_27342 = ~n_27332 & ~n_27341;
assign n_27343 = ~n_27331 & ~n_27342;
assign n_27344 = ~n_27330 & ~n_27343;
assign n_27345 = ~n_27329 & ~n_27344;
assign n_27346 = ~n_27328 & ~n_27345;
assign n_27347 = ~n_27327 & ~n_27346;
assign n_27348 = ~n_27326 & ~n_27347;
assign n_27349 = ~n_27325 & ~n_27348;
assign n_27350 = ~n_27324 & ~n_27349;
assign n_27351 = ~n_27323 & ~n_27350;
assign n_27352 = ~n_27322 & ~n_27351;
assign n_27353 = ~n_27321 & ~n_27352;
assign n_27354 = ~n_27320 & ~n_27353;
assign n_27355 = ~n_27319 & ~n_27354;
assign n_27356 = ~n_27318 & ~n_27355;
assign n_27357 = ~n_27317 & ~n_27356;
assign n_27358 = ~n_27316 & ~n_27357;
assign n_27359 = ~n_27315 & ~n_27358;
assign n_27360 = ~n_27314 & ~n_27359;
assign n_27361 = ~n_27313 & ~n_27360;
assign n_27362 = ~n_27312 & ~n_27361;
assign n_27363 = ~n_27311 & ~n_27362;
assign n_27364 = ~n_27310 & ~n_27363;
assign n_27365 = ~n_27309 & ~n_27364;
assign n_27366 = ~n_27308 & ~n_27365;
assign n_27367 = ~n_27307 & ~n_27366;
assign n_27368 = ~n_27306 & ~n_27367;
assign n_27369 = ~n_27305 & ~n_27368;
assign n_27370 = ~n_27304 & ~n_27369;
assign n_27371 = ~n_27303 & ~n_27370;
assign n_27372 = ~n_27302 & ~n_27371;
assign n_27373 = ~n_27301 & ~n_27372;
assign n_27374 = ~n_27300 & ~n_27373;
assign n_27375 = ~n_27299 & ~n_27374;
assign n_27376 = ~n_27298 & ~n_27375;
assign n_27377 = ~n_27297 & ~n_27376;
assign n_27378 = ~n_27296 & ~n_27377;
assign n_27379 = ~n_27295 & ~n_27378;
assign n_27380 = ~n_27294 & ~n_27379;
assign n_27381 = ~n_27293 & ~n_27380;
assign n_27382 = ~n_27292 & ~n_27381;
assign n_27383 = ~n_27291 & ~n_27382;
assign n_27384 = ~n_27290 & ~n_27383;
assign n_27385 = ~n_27289 & ~n_27384;
assign n_27386 = ~n_27288 & ~n_27385;
assign n_27387 = ~n_27287 & ~n_27386;
assign n_27388 = ~n_27286 & ~n_27387;
assign n_27389 = ~n_27285 & ~n_27388;
assign n_27390 = ~n_27284 & ~n_27389;
assign n_27391 = ~n_27283 & ~n_27390;
assign n_27392 = ~n_27282 & ~n_27391;
assign n_27393 = ~n_27281 & ~n_27392;
assign n_27394 = ~n_27280 & ~n_27393;
assign n_27395 = ~n_27279 & ~n_27394;
assign n_27396 = ~n_27278 & ~n_27395;
assign n_27397 = ~n_27277 & ~n_27396;
assign n_27398 = ~n_27276 & ~n_27397;
assign n_27399 = ~n_27275 & ~n_27398;
assign n_27400 = ~n_27399 &  n_19945;
assign n_27401 =  n_27274 &  n_27400;
assign n_27402 =  x_37 &  n_27273;
assign n_27403 = ~x_38 &  n_27402;
assign n_27404 =  n_3664 &  n_27403;
assign n_27405 =  n_27254 &  n_27404;
assign n_27406 =  n_389 &  n_7;
assign n_27407 =  n_12420 &  n_27406;
assign n_27408 = ~n_27399 &  n_27407;
assign n_27409 = ~n_27405 & ~n_27408;
assign n_27410 = ~n_27401 &  n_27409;
assign n_27411 = ~n_27399 &  n_27403;
assign n_27412 =  n_12420 &  n_27411;
assign n_27413 =  x_38 &  n_27266;
assign n_27414 =  n_3664 &  n_27413;
assign n_27415 =  n_27254 &  n_27414;
assign n_27416 =  x_38 &  n_27274;
assign n_27417 =  n_8818 &  n_27416;
assign n_27418 = ~n_27254 &  n_27417;
assign n_27419 = ~n_27415 & ~n_27418;
assign n_27420 = ~n_27412 &  n_27419;
assign n_27421 =  n_27410 &  n_27420;
assign n_27422 = ~x_36 &  x_37;
assign n_27423 =  n_27256 &  n_27422;
assign n_27424 = ~x_38 &  n_27423;
assign n_27425 =  n_8818 &  n_27424;
assign n_27426 =  n_27254 &  n_27425;
assign n_27427 = ~x_336 &  x_1424;
assign n_27428 =  x_337 & ~x_1425;
assign n_27429 = ~x_337 &  x_1425;
assign n_27430 =  x_338 & ~x_1426;
assign n_27431 = ~x_338 &  x_1426;
assign n_27432 =  x_339 & ~x_1427;
assign n_27433 = ~x_339 &  x_1427;
assign n_27434 =  x_340 & ~x_1428;
assign n_27435 = ~x_340 &  x_1428;
assign n_27436 =  x_341 & ~x_1429;
assign n_27437 = ~x_341 &  x_1429;
assign n_27438 =  x_342 & ~x_1430;
assign n_27439 = ~x_342 &  x_1430;
assign n_27440 =  x_343 & ~x_1431;
assign n_27441 = ~x_343 &  x_1431;
assign n_27442 =  x_344 & ~x_1432;
assign n_27443 = ~x_344 &  x_1432;
assign n_27444 =  x_345 & ~x_1433;
assign n_27445 = ~x_345 &  x_1433;
assign n_27446 =  x_346 & ~x_1434;
assign n_27447 = ~x_346 &  x_1434;
assign n_27448 =  x_347 & ~x_1435;
assign n_27449 = ~x_347 &  x_1435;
assign n_27450 =  x_348 & ~x_1436;
assign n_27451 = ~x_348 &  x_1436;
assign n_27452 =  x_349 & ~x_1437;
assign n_27453 = ~x_349 &  x_1437;
assign n_27454 =  x_350 & ~x_1438;
assign n_27455 = ~x_350 &  x_1438;
assign n_27456 =  x_351 & ~x_1439;
assign n_27457 = ~x_351 &  x_1439;
assign n_27458 =  x_352 & ~x_1440;
assign n_27459 = ~x_352 &  x_1440;
assign n_27460 =  x_353 & ~x_1441;
assign n_27461 = ~x_353 &  x_1441;
assign n_27462 =  x_354 & ~x_1442;
assign n_27463 = ~x_354 &  x_1442;
assign n_27464 =  x_355 & ~x_1443;
assign n_27465 = ~x_355 &  x_1443;
assign n_27466 =  x_356 & ~x_1444;
assign n_27467 = ~x_356 &  x_1444;
assign n_27468 =  x_357 & ~x_1445;
assign n_27469 = ~x_357 &  x_1445;
assign n_27470 =  x_358 & ~x_1446;
assign n_27471 = ~x_358 &  x_1446;
assign n_27472 =  x_359 & ~x_1447;
assign n_27473 = ~x_359 &  x_1447;
assign n_27474 =  x_361 & ~x_1449;
assign n_27475 = ~x_362 &  x_1450;
assign n_27476 = ~n_27474 &  n_27475;
assign n_27477 = ~x_361 &  x_1449;
assign n_27478 = ~x_360 &  x_1448;
assign n_27479 = ~n_27477 & ~n_27478;
assign n_27480 = ~n_27476 &  n_27479;
assign n_27481 =  x_360 & ~x_1448;
assign n_27482 = ~n_27480 & ~n_27481;
assign n_27483 = ~n_27473 & ~n_27482;
assign n_27484 = ~n_27472 & ~n_27483;
assign n_27485 = ~n_27471 & ~n_27484;
assign n_27486 = ~n_27470 & ~n_27485;
assign n_27487 = ~n_27469 & ~n_27486;
assign n_27488 = ~n_27468 & ~n_27487;
assign n_27489 = ~n_27467 & ~n_27488;
assign n_27490 = ~n_27466 & ~n_27489;
assign n_27491 = ~n_27465 & ~n_27490;
assign n_27492 = ~n_27464 & ~n_27491;
assign n_27493 = ~n_27463 & ~n_27492;
assign n_27494 = ~n_27462 & ~n_27493;
assign n_27495 = ~n_27461 & ~n_27494;
assign n_27496 = ~n_27460 & ~n_27495;
assign n_27497 = ~n_27459 & ~n_27496;
assign n_27498 = ~n_27458 & ~n_27497;
assign n_27499 = ~n_27457 & ~n_27498;
assign n_27500 = ~n_27456 & ~n_27499;
assign n_27501 = ~n_27455 & ~n_27500;
assign n_27502 = ~n_27454 & ~n_27501;
assign n_27503 = ~n_27453 & ~n_27502;
assign n_27504 = ~n_27452 & ~n_27503;
assign n_27505 = ~n_27451 & ~n_27504;
assign n_27506 = ~n_27450 & ~n_27505;
assign n_27507 = ~n_27449 & ~n_27506;
assign n_27508 = ~n_27448 & ~n_27507;
assign n_27509 = ~n_27447 & ~n_27508;
assign n_27510 = ~n_27446 & ~n_27509;
assign n_27511 = ~n_27445 & ~n_27510;
assign n_27512 = ~n_27444 & ~n_27511;
assign n_27513 = ~n_27443 & ~n_27512;
assign n_27514 = ~n_27442 & ~n_27513;
assign n_27515 = ~n_27441 & ~n_27514;
assign n_27516 = ~n_27440 & ~n_27515;
assign n_27517 = ~n_27439 & ~n_27516;
assign n_27518 = ~n_27438 & ~n_27517;
assign n_27519 = ~n_27437 & ~n_27518;
assign n_27520 = ~n_27436 & ~n_27519;
assign n_27521 = ~n_27435 & ~n_27520;
assign n_27522 = ~n_27434 & ~n_27521;
assign n_27523 = ~n_27433 & ~n_27522;
assign n_27524 = ~n_27432 & ~n_27523;
assign n_27525 = ~n_27431 & ~n_27524;
assign n_27526 = ~n_27430 & ~n_27525;
assign n_27527 = ~n_27429 & ~n_27526;
assign n_27528 = ~n_27428 & ~n_27527;
assign n_27529 = ~n_27427 & ~n_27528;
assign n_27530 =  x_336 & ~x_1424;
assign n_27531 =  x_335 & ~x_1423;
assign n_27532 = ~n_27530 & ~n_27531;
assign n_27533 = ~n_27529 &  n_27532;
assign n_27534 = ~x_334 &  x_1422;
assign n_27535 = ~x_335 &  x_1423;
assign n_27536 = ~n_27534 & ~n_27535;
assign n_27537 = ~n_27533 &  n_27536;
assign n_27538 =  x_334 & ~x_1422;
assign n_27539 =  x_333 & ~x_1421;
assign n_27540 = ~n_27538 & ~n_27539;
assign n_27541 = ~n_27537 &  n_27540;
assign n_27542 = ~x_332 &  x_1420;
assign n_27543 = ~x_333 &  x_1421;
assign n_27544 = ~n_27542 & ~n_27543;
assign n_27545 = ~n_27541 &  n_27544;
assign n_27546 =  x_332 & ~x_1420;
assign n_27547 = ~x_331 &  x_1419;
assign n_27548 = ~n_27546 & ~n_27547;
assign n_27549 = ~n_27545 &  n_27548;
assign n_27550 =  n_24801 &  n_1179;
assign n_27551 =  x_331 & ~x_1419;
assign n_27552 =  n_27550 & ~n_27551;
assign n_27553 = ~n_27549 &  n_27552;
assign n_27554 = ~x_1982 & ~x_1983;
assign n_27555 = ~x_1984 & ~x_1985;
assign n_27556 =  n_27554 &  n_27555;
assign n_27557 = ~x_1978 & ~x_1979;
assign n_27558 = ~x_1980 & ~x_1981;
assign n_27559 =  n_27557 &  n_27558;
assign n_27560 =  n_27556 &  n_27559;
assign n_27561 = ~x_1990 & ~x_1991;
assign n_27562 = ~x_1992 &  n_27561;
assign n_27563 = ~x_1986 & ~x_1987;
assign n_27564 = ~x_1988 & ~x_1989;
assign n_27565 =  n_27563 &  n_27564;
assign n_27566 =  n_27562 &  n_27565;
assign n_27567 =  n_27560 &  n_27566;
assign n_27568 = ~x_1964 & ~x_1965;
assign n_27569 = ~x_1966 & ~x_1967;
assign n_27570 = ~x_1968 & ~x_1969;
assign n_27571 =  n_27569 &  n_27570;
assign n_27572 =  n_27568 &  n_27571;
assign n_27573 = ~x_1974 & ~x_1975;
assign n_27574 = ~x_1976 & ~x_1977;
assign n_27575 =  n_27573 &  n_27574;
assign n_27576 = ~x_1970 & ~x_1971;
assign n_27577 = ~x_1972 & ~x_1973;
assign n_27578 =  n_27576 &  n_27577;
assign n_27579 =  n_27575 &  n_27578;
assign n_27580 =  n_27572 &  n_27579;
assign n_27581 =  n_27567 &  n_27580;
assign n_27582 = ~x_1963 & ~n_27581;
assign n_27583 =  n_982 &  n_18445;
assign n_27584 = ~n_27582 &  n_27583;
assign n_27585 = ~x_39 &  n_983;
assign n_27586 = ~x_40 &  n_27585;
assign n_27587 =  n_4992 &  n_27586;
assign n_27588 =  n_3469 &  n_18439;
assign n_27589 = ~n_27588 & ~n_984;
assign n_27590 = ~n_27587 &  n_27589;
assign n_27591 = ~n_27584 &  n_27590;
assign n_27592 =  n_980 &  n_6527;
assign n_27593 = ~x_39 &  n_27267;
assign n_27594 =  n_27593 &  n_12614;
assign n_27595 = ~n_27592 & ~n_27594;
assign n_27596 =  n_1906 &  n_27416;
assign n_27597 = ~n_192 & ~n_27596;
assign n_27598 =  n_1315 &  n_27593;
assign n_27599 =  x_38 &  n_27423;
assign n_27600 =  x_39 &  n_1706;
assign n_27601 =  n_27599 &  n_27600;
assign n_27602 =  x_40 &  n_27601;
assign n_27603 = ~n_27598 & ~n_27602;
assign n_27604 =  n_27597 &  n_27603;
assign n_27605 =  n_27595 &  n_27604;
assign n_27606 =  n_27591 &  n_27605;
assign n_27607 = ~x_1151 & ~x_1152;
assign n_27608 = ~x_1153 & ~x_1154;
assign n_27609 =  n_27607 &  n_27608;
assign n_27610 = ~x_1147 & ~x_1148;
assign n_27611 = ~x_1149 & ~x_1150;
assign n_27612 =  n_27610 &  n_27611;
assign n_27613 =  n_27609 &  n_27612;
assign n_27614 = ~x_1159 & ~x_1160;
assign n_27615 = ~x_1161 & ~x_1162;
assign n_27616 =  n_27614 &  n_27615;
assign n_27617 = ~x_1155 & ~x_1156;
assign n_27618 = ~x_1157 & ~x_1158;
assign n_27619 =  n_27617 &  n_27618;
assign n_27620 =  n_27616 &  n_27619;
assign n_27621 =  n_27613 &  n_27620;
assign n_27622 = ~x_1135 & ~x_1136;
assign n_27623 = ~x_1137 & ~x_1138;
assign n_27624 =  n_27622 &  n_27623;
assign n_27625 = ~x_1131 & ~x_1132;
assign n_27626 = ~x_1133 & ~x_1134;
assign n_27627 =  n_27625 &  n_27626;
assign n_27628 =  n_27624 &  n_27627;
assign n_27629 = ~x_1143 & ~x_1144;
assign n_27630 = ~x_1145 & ~x_1146;
assign n_27631 =  n_27629 &  n_27630;
assign n_27632 = ~x_1139 & ~x_1140;
assign n_27633 = ~x_1141 & ~x_1142;
assign n_27634 =  n_27632 &  n_27633;
assign n_27635 =  n_27631 &  n_27634;
assign n_27636 =  n_27628 &  n_27635;
assign n_27637 =  n_27621 &  n_27636;
assign n_27638 =  n_2101 & ~n_27637;
assign n_27639 =  n_3664 &  n_27638;
assign n_27640 = ~x_350 & ~x_351;
assign n_27641 = ~x_352 & ~x_353;
assign n_27642 =  n_27640 &  n_27641;
assign n_27643 = ~x_346 & ~x_347;
assign n_27644 = ~x_348 & ~x_349;
assign n_27645 =  n_27643 &  n_27644;
assign n_27646 =  n_27642 &  n_27645;
assign n_27647 = ~x_358 & ~x_359;
assign n_27648 = ~x_360 &  n_27647;
assign n_27649 = ~x_354 & ~x_355;
assign n_27650 = ~x_356 & ~x_357;
assign n_27651 =  n_27649 &  n_27650;
assign n_27652 =  n_27648 &  n_27651;
assign n_27653 =  n_27646 &  n_27652;
assign n_27654 = ~x_332 & ~x_333;
assign n_27655 = ~x_334 & ~x_335;
assign n_27656 = ~x_336 & ~x_337;
assign n_27657 =  n_27655 &  n_27656;
assign n_27658 =  n_27654 &  n_27657;
assign n_27659 = ~x_342 & ~x_343;
assign n_27660 = ~x_344 & ~x_345;
assign n_27661 =  n_27659 &  n_27660;
assign n_27662 = ~x_338 & ~x_339;
assign n_27663 = ~x_340 & ~x_341;
assign n_27664 =  n_27662 &  n_27663;
assign n_27665 =  n_27661 &  n_27664;
assign n_27666 =  n_27658 &  n_27665;
assign n_27667 =  n_27653 &  n_27666;
assign n_27668 = ~x_361 &  n_27667;
assign n_27669 = ~x_331 & ~n_27668;
assign n_27670 =  n_12420 &  n_2101;
assign n_27671 = ~n_27669 &  n_27670;
assign n_27672 = ~n_27639 & ~n_27671;
assign n_27673 = ~x_1087 & ~x_1088;
assign n_27674 = ~x_1089 & ~x_1090;
assign n_27675 =  n_27673 &  n_27674;
assign n_27676 = ~x_1083 & ~x_1084;
assign n_27677 = ~x_1085 & ~x_1086;
assign n_27678 =  n_27676 &  n_27677;
assign n_27679 =  n_27675 &  n_27678;
assign n_27680 = ~x_1095 & ~x_1096;
assign n_27681 = ~x_1097 & ~x_1098;
assign n_27682 =  n_27680 &  n_27681;
assign n_27683 = ~x_1091 & ~x_1092;
assign n_27684 = ~x_1093 & ~x_1094;
assign n_27685 =  n_27683 &  n_27684;
assign n_27686 =  n_27682 &  n_27685;
assign n_27687 =  n_27679 &  n_27686;
assign n_27688 = ~x_1071 & ~x_1072;
assign n_27689 = ~x_1073 & ~x_1074;
assign n_27690 =  n_27688 &  n_27689;
assign n_27691 = ~x_1067 & ~x_1068;
assign n_27692 = ~x_1069 & ~x_1070;
assign n_27693 =  n_27691 &  n_27692;
assign n_27694 =  n_27690 &  n_27693;
assign n_27695 = ~x_1079 & ~x_1080;
assign n_27696 = ~x_1081 & ~x_1082;
assign n_27697 =  n_27695 &  n_27696;
assign n_27698 = ~x_1075 & ~x_1076;
assign n_27699 = ~x_1077 & ~x_1078;
assign n_27700 =  n_27698 &  n_27699;
assign n_27701 =  n_27697 &  n_27700;
assign n_27702 =  n_27694 &  n_27701;
assign n_27703 =  n_27687 &  n_27702;
assign n_27704 =  n_191 & ~n_27703;
assign n_27705 =  n_1707 &  n_27704;
assign n_27706 =  n_3 &  n_3275;
assign n_27707 = ~n_4446 & ~n_27706;
assign n_27708 =  n_10318 &  n_8803;
assign n_27709 = ~n_19946 & ~n_27708;
assign n_27710 =  n_27707 &  n_27709;
assign n_27711 =  n_6533 &  n_27416;
assign n_27712 = ~n_23504 & ~n_27711;
assign n_27713 =  n_27710 &  n_27712;
assign n_27714 = ~n_27705 &  n_27713;
assign n_27715 =  n_27672 &  n_27714;
assign n_27716 =  n_27606 &  n_27715;
assign n_27717 = ~x_1438 & ~x_1439;
assign n_27718 = ~x_1440 & ~x_1441;
assign n_27719 =  n_27717 &  n_27718;
assign n_27720 = ~x_1434 & ~x_1435;
assign n_27721 = ~x_1436 & ~x_1437;
assign n_27722 =  n_27720 &  n_27721;
assign n_27723 =  n_27719 &  n_27722;
assign n_27724 = ~x_1446 & ~x_1447;
assign n_27725 = ~x_1448 &  n_27724;
assign n_27726 = ~x_1442 & ~x_1443;
assign n_27727 = ~x_1444 & ~x_1445;
assign n_27728 =  n_27726 &  n_27727;
assign n_27729 =  n_27725 &  n_27728;
assign n_27730 =  n_27723 &  n_27729;
assign n_27731 = ~x_1420 & ~x_1421;
assign n_27732 = ~x_1422 & ~x_1423;
assign n_27733 = ~x_1424 & ~x_1425;
assign n_27734 =  n_27732 &  n_27733;
assign n_27735 =  n_27731 &  n_27734;
assign n_27736 = ~x_1430 & ~x_1431;
assign n_27737 = ~x_1432 & ~x_1433;
assign n_27738 =  n_27736 &  n_27737;
assign n_27739 = ~x_1426 & ~x_1427;
assign n_27740 = ~x_1428 & ~x_1429;
assign n_27741 =  n_27739 &  n_27740;
assign n_27742 =  n_27738 &  n_27741;
assign n_27743 =  n_27735 &  n_27742;
assign n_27744 =  n_27730 &  n_27743;
assign n_27745 = ~x_1449 &  n_27744;
assign n_27746 = ~x_1419 & ~n_27745;
assign n_27747 =  n_1903 & ~n_27746;
assign n_27748 =  n_3664 &  n_389;
assign n_27749 =  n_27747 &  n_27748;
assign n_27750 = ~x_511 & ~x_512;
assign n_27751 = ~x_513 & ~x_514;
assign n_27752 =  n_27750 &  n_27751;
assign n_27753 = ~x_507 & ~x_508;
assign n_27754 = ~x_509 & ~x_510;
assign n_27755 =  n_27753 &  n_27754;
assign n_27756 =  n_27752 &  n_27755;
assign n_27757 = ~x_519 & ~x_520;
assign n_27758 = ~x_521 & ~x_522;
assign n_27759 =  n_27757 &  n_27758;
assign n_27760 = ~x_515 & ~x_516;
assign n_27761 = ~x_517 & ~x_518;
assign n_27762 =  n_27760 &  n_27761;
assign n_27763 =  n_27759 &  n_27762;
assign n_27764 =  n_27756 &  n_27763;
assign n_27765 = ~x_495 & ~x_496;
assign n_27766 = ~x_497 & ~x_498;
assign n_27767 =  n_27765 &  n_27766;
assign n_27768 = ~x_491 & ~x_492;
assign n_27769 = ~x_493 & ~x_494;
assign n_27770 =  n_27768 &  n_27769;
assign n_27771 =  n_27767 &  n_27770;
assign n_27772 = ~x_503 & ~x_504;
assign n_27773 = ~x_505 & ~x_506;
assign n_27774 =  n_27772 &  n_27773;
assign n_27775 = ~x_499 & ~x_500;
assign n_27776 = ~x_501 & ~x_502;
assign n_27777 =  n_27775 &  n_27776;
assign n_27778 =  n_27774 &  n_27777;
assign n_27779 =  n_27771 &  n_27778;
assign n_27780 =  n_27764 &  n_27779;
assign n_27781 =  n_2 &  n_18433;
assign n_27782 =  n_27780 &  n_27781;
assign n_27783 = ~x_1118 & ~x_1119;
assign n_27784 = ~x_1120 & ~x_1121;
assign n_27785 =  n_27783 &  n_27784;
assign n_27786 = ~x_1114 & ~x_1115;
assign n_27787 = ~x_1116 & ~x_1117;
assign n_27788 =  n_27786 &  n_27787;
assign n_27789 =  n_27785 &  n_27788;
assign n_27790 = ~x_1126 & ~x_1127;
assign n_27791 = ~x_1128 &  n_27790;
assign n_27792 = ~x_1122 & ~x_1123;
assign n_27793 = ~x_1124 & ~x_1125;
assign n_27794 =  n_27792 &  n_27793;
assign n_27795 =  n_27791 &  n_27794;
assign n_27796 =  n_27789 &  n_27795;
assign n_27797 = ~x_1100 & ~x_1101;
assign n_27798 = ~x_1102 & ~x_1103;
assign n_27799 = ~x_1104 & ~x_1105;
assign n_27800 =  n_27798 &  n_27799;
assign n_27801 =  n_27797 &  n_27800;
assign n_27802 = ~x_1110 & ~x_1111;
assign n_27803 = ~x_1112 & ~x_1113;
assign n_27804 =  n_27802 &  n_27803;
assign n_27805 = ~x_1106 & ~x_1107;
assign n_27806 = ~x_1108 & ~x_1109;
assign n_27807 =  n_27805 &  n_27806;
assign n_27808 =  n_27804 &  n_27807;
assign n_27809 =  n_27801 &  n_27808;
assign n_27810 =  n_27796 &  n_27809;
assign n_27811 = ~x_1099 & ~n_27810;
assign n_27812 = ~x_33 & ~n_27811;
assign n_27813 =  n_2886 &  n_3859;
assign n_27814 =  n_12614 &  n_27813;
assign n_27815 = ~x_34 &  x_35;
assign n_27816 =  n_27814 &  n_27815;
assign n_27817 =  n_27812 &  n_27816;
assign n_27818 = ~n_27782 & ~n_27817;
assign n_27819 = ~n_27749 &  n_27818;
assign n_27820 =  n_783 &  n_4;
assign n_27821 =  n_1903 &  n_27746;
assign n_27822 =  n_27820 &  n_27821;
assign n_27823 =  n_2101 &  n_27637;
assign n_27824 =  n_980 &  n_27823;
assign n_27825 =  n_12420 &  n_191;
assign n_27826 = ~n_27669 &  n_27825;
assign n_27827 = ~n_27824 & ~n_27826;
assign n_27828 = ~n_27822 &  n_27827;
assign n_27829 =  n_27819 &  n_27828;
assign n_27830 =  n_27716 &  n_27829;
assign n_27831 = ~x_1450 &  n_27745;
assign n_27832 = ~x_1419 & ~n_27831;
assign n_27833 =  n_1903 & ~n_27832;
assign n_27834 =  n_24413 &  n_27833;
assign n_27835 =  n_4993 &  n_1904;
assign n_27836 =  n_27780 &  n_27835;
assign n_27837 = ~n_27834 & ~n_27836;
assign n_27838 =  x_42 &  n_20718;
assign n_27839 =  n_3 &  n_12226;
assign n_27840 =  n_3663 &  n_983;
assign n_27841 =  x_42 &  n_27840;
assign n_27842 = ~n_27839 & ~n_27841;
assign n_27843 = ~n_27838 &  n_27842;
assign n_27844 = ~x_2207 & ~x_2208;
assign n_27845 = ~x_2209 & ~x_2210;
assign n_27846 =  n_27844 &  n_27845;
assign n_27847 = ~x_2203 & ~x_2204;
assign n_27848 = ~x_2205 & ~x_2206;
assign n_27849 =  n_27847 &  n_27848;
assign n_27850 =  n_27846 &  n_27849;
assign n_27851 = ~x_2215 & ~x_2216;
assign n_27852 = ~x_2217 & ~x_2218;
assign n_27853 =  n_27851 &  n_27852;
assign n_27854 = ~x_2211 & ~x_2212;
assign n_27855 = ~x_2213 & ~x_2214;
assign n_27856 =  n_27854 &  n_27855;
assign n_27857 =  n_27853 &  n_27856;
assign n_27858 =  n_27850 &  n_27857;
assign n_27859 = ~x_2191 & ~x_2192;
assign n_27860 = ~x_2193 & ~x_2194;
assign n_27861 =  n_27859 &  n_27860;
assign n_27862 = ~x_2187 & ~x_2188;
assign n_27863 = ~x_2189 & ~x_2190;
assign n_27864 =  n_27862 &  n_27863;
assign n_27865 =  n_27861 &  n_27864;
assign n_27866 = ~x_2199 & ~x_2200;
assign n_27867 = ~x_2201 & ~x_2202;
assign n_27868 =  n_27866 &  n_27867;
assign n_27869 = ~x_2195 & ~x_2196;
assign n_27870 = ~x_2197 & ~x_2198;
assign n_27871 =  n_27869 &  n_27870;
assign n_27872 =  n_27868 &  n_27871;
assign n_27873 =  n_27865 &  n_27872;
assign n_27874 =  n_27858 &  n_27873;
assign n_27875 =  n_3469 &  n_983;
assign n_27876 = ~n_27874 &  n_27875;
assign n_27877 =  n_587 &  n_4057;
assign n_27878 = ~x_831 & ~x_832;
assign n_27879 = ~x_833 & ~x_834;
assign n_27880 =  n_27878 &  n_27879;
assign n_27881 = ~x_827 & ~x_828;
assign n_27882 = ~x_829 & ~x_830;
assign n_27883 =  n_27881 &  n_27882;
assign n_27884 =  n_27880 &  n_27883;
assign n_27885 = ~x_839 & ~x_840;
assign n_27886 = ~x_841 & ~x_842;
assign n_27887 =  n_27885 &  n_27886;
assign n_27888 = ~x_835 & ~x_836;
assign n_27889 = ~x_837 & ~x_838;
assign n_27890 =  n_27888 &  n_27889;
assign n_27891 =  n_27887 &  n_27890;
assign n_27892 =  n_27884 &  n_27891;
assign n_27893 = ~x_815 & ~x_816;
assign n_27894 = ~x_817 & ~x_818;
assign n_27895 =  n_27893 &  n_27894;
assign n_27896 = ~x_811 & ~x_812;
assign n_27897 = ~x_813 & ~x_814;
assign n_27898 =  n_27896 &  n_27897;
assign n_27899 =  n_27895 &  n_27898;
assign n_27900 = ~x_823 & ~x_824;
assign n_27901 = ~x_825 & ~x_826;
assign n_27902 =  n_27900 &  n_27901;
assign n_27903 = ~x_819 & ~x_820;
assign n_27904 = ~x_821 & ~x_822;
assign n_27905 =  n_27903 &  n_27904;
assign n_27906 =  n_27902 &  n_27905;
assign n_27907 =  n_27899 &  n_27906;
assign n_27908 =  n_27892 &  n_27907;
assign n_27909 =  n_27877 & ~n_27908;
assign n_27910 = ~n_27876 & ~n_27909;
assign n_27911 =  n_27413 &  n_1707;
assign n_27912 =  x_42 &  n_23894;
assign n_27913 = ~n_27911 & ~n_27912;
assign n_27914 =  n_27910 &  n_27913;
assign n_27915 =  n_27843 &  n_27914;
assign n_27916 =  n_980 &  n_18439;
assign n_27917 =  x_1449 &  x_1450;
assign n_27918 =  n_27744 & ~n_27917;
assign n_27919 = ~x_1419 & ~n_27918;
assign n_27920 =  n_27916 & ~n_27919;
assign n_27921 = ~n_8808 & ~n_27920;
assign n_27922 =  n_27915 &  n_27921;
assign n_27923 = ~n_2102 & ~n_13860;
assign n_27924 =  n_782 &  n_983;
assign n_27925 =  n_4992 &  n_27924;
assign n_27926 = ~n_3863 & ~n_12033;
assign n_27927 = ~n_6529 &  n_27926;
assign n_27928 = ~n_27925 &  n_27927;
assign n_27929 =  n_27923 &  n_27928;
assign n_27930 =  x_34 & ~x_35;
assign n_27931 =  n_3859 &  n_27930;
assign n_27932 =  n_6530 &  n_27931;
assign n_27933 =  n_27812 &  n_27932;
assign n_27934 =  n_2 &  n_4251;
assign n_27935 = ~n_27933 & ~n_27934;
assign n_27936 =  n_27929 &  n_27935;
assign n_27937 =  n_27922 &  n_27936;
assign n_27938 =  n_27837 &  n_27937;
assign n_27939 =  n_27830 &  n_27938;
assign n_27940 = ~x_1503 & ~x_1504;
assign n_27941 = ~x_1505 & ~x_1506;
assign n_27942 =  n_27940 &  n_27941;
assign n_27943 = ~x_1499 & ~x_1500;
assign n_27944 = ~x_1501 & ~x_1502;
assign n_27945 =  n_27943 &  n_27944;
assign n_27946 =  n_27942 &  n_27945;
assign n_27947 = ~x_1511 & ~x_1512;
assign n_27948 = ~x_1513 & ~x_1514;
assign n_27949 =  n_27947 &  n_27948;
assign n_27950 = ~x_1507 & ~x_1508;
assign n_27951 = ~x_1509 & ~x_1510;
assign n_27952 =  n_27950 &  n_27951;
assign n_27953 =  n_27949 &  n_27952;
assign n_27954 =  n_27946 &  n_27953;
assign n_27955 = ~x_1487 & ~x_1488;
assign n_27956 = ~x_1489 & ~x_1490;
assign n_27957 =  n_27955 &  n_27956;
assign n_27958 = ~x_1483 & ~x_1484;
assign n_27959 = ~x_1485 & ~x_1486;
assign n_27960 =  n_27958 &  n_27959;
assign n_27961 =  n_27957 &  n_27960;
assign n_27962 = ~x_1495 & ~x_1496;
assign n_27963 = ~x_1497 & ~x_1498;
assign n_27964 =  n_27962 &  n_27963;
assign n_27965 = ~x_1491 & ~x_1492;
assign n_27966 = ~x_1493 & ~x_1494;
assign n_27967 =  n_27965 &  n_27966;
assign n_27968 =  n_27964 &  n_27967;
assign n_27969 =  n_27961 &  n_27968;
assign n_27970 =  n_27954 &  n_27969;
assign n_27971 =  n_1709 &  n_27970;
assign n_27972 =  n_8060 &  n_27971;
assign n_27973 = ~x_1099 &  n_5;
assign n_27974 =  x_1129 &  x_1130;
assign n_27975 =  n_27810 & ~n_27974;
assign n_27976 =  n_27973 & ~n_27975;
assign n_27977 =  n_188 &  n_8255;
assign n_27978 =  n_27976 &  n_27977;
assign n_27979 = ~n_27972 & ~n_27978;
assign n_27980 = ~x_767 & ~x_768;
assign n_27981 = ~x_769 & ~x_770;
assign n_27982 =  n_27980 &  n_27981;
assign n_27983 = ~x_763 & ~x_764;
assign n_27984 = ~x_765 & ~x_766;
assign n_27985 =  n_27983 &  n_27984;
assign n_27986 =  n_27982 &  n_27985;
assign n_27987 = ~x_775 & ~x_776;
assign n_27988 = ~x_777 & ~x_778;
assign n_27989 =  n_27987 &  n_27988;
assign n_27990 = ~x_771 & ~x_772;
assign n_27991 = ~x_773 & ~x_774;
assign n_27992 =  n_27990 &  n_27991;
assign n_27993 =  n_27989 &  n_27992;
assign n_27994 =  n_27986 &  n_27993;
assign n_27995 = ~x_751 & ~x_752;
assign n_27996 = ~x_753 & ~x_754;
assign n_27997 =  n_27995 &  n_27996;
assign n_27998 = ~x_747 & ~x_748;
assign n_27999 = ~x_749 & ~x_750;
assign n_28000 =  n_27998 &  n_27999;
assign n_28001 =  n_27997 &  n_28000;
assign n_28002 = ~x_759 & ~x_760;
assign n_28003 = ~x_761 & ~x_762;
assign n_28004 =  n_28002 &  n_28003;
assign n_28005 = ~x_755 & ~x_756;
assign n_28006 = ~x_757 & ~x_758;
assign n_28007 =  n_28005 &  n_28006;
assign n_28008 =  n_28004 &  n_28007;
assign n_28009 =  n_28001 &  n_28008;
assign n_28010 =  n_7 &  n_28009;
assign n_28011 =  n_27994 &  n_28010;
assign n_28012 =  n_10318 &  n_2302;
assign n_28013 =  n_28011 &  n_28012;
assign n_28014 = ~x_1963 &  n_387;
assign n_28015 =  x_1993 &  x_1994;
assign n_28016 =  n_27581 & ~n_28015;
assign n_28017 =  n_28014 & ~n_28016;
assign n_28018 =  n_3858 &  n_13005;
assign n_28019 =  n_28017 &  n_28018;
assign n_28020 = ~n_28013 & ~n_28019;
assign n_28021 =  n_27979 &  n_28020;
assign n_28022 =  n_2100 &  n_24801;
assign n_28023 =  n_1903 &  n_27832;
assign n_28024 =  n_28022 &  n_28023;
assign n_28025 =  n_28021 & ~n_28024;
assign n_28026 =  n_980 &  n_27638;
assign n_28027 =  n_13012 &  n_8802;
assign n_28028 = ~x_362 &  n_27668;
assign n_28029 = ~x_331 & ~n_28028;
assign n_28030 =  n_28027 & ~n_28029;
assign n_28031 = ~n_28026 & ~n_28030;
assign n_28032 =  x_361 &  x_362;
assign n_28033 =  n_27667 & ~n_28032;
assign n_28034 = ~x_331 & ~n_28033;
assign n_28035 =  n_12614 &  n_10518;
assign n_28036 =  n_28034 &  n_28035;
assign n_28037 = ~x_331 & ~n_27667;
assign n_28038 =  n_980 &  n_1179;
assign n_28039 = ~n_28037 &  n_28038;
assign n_28040 =  n_3664 &  n_27823;
assign n_28041 = ~n_1706 &  n_1180;
assign n_28042 = ~n_28040 & ~n_28041;
assign n_28043 = ~n_28039 &  n_28042;
assign n_28044 = ~n_28036 &  n_28043;
assign n_28045 =  n_28031 &  n_28044;
assign n_28046 =  n_28025 &  n_28045;
assign n_28047 =  n_1315 &  n_2303;
assign n_28048 = ~x_2431 & ~x_2432;
assign n_28049 = ~x_2433 & ~x_2434;
assign n_28050 =  n_28048 &  n_28049;
assign n_28051 = ~x_2427 & ~x_2428;
assign n_28052 = ~x_2429 & ~x_2430;
assign n_28053 =  n_28051 &  n_28052;
assign n_28054 =  n_28050 &  n_28053;
assign n_28055 = ~x_2439 & ~x_2440;
assign n_28056 = ~x_2441 & ~x_2442;
assign n_28057 =  n_28055 &  n_28056;
assign n_28058 = ~x_2435 & ~x_2436;
assign n_28059 = ~x_2437 & ~x_2438;
assign n_28060 =  n_28058 &  n_28059;
assign n_28061 =  n_28057 &  n_28060;
assign n_28062 =  n_28054 &  n_28061;
assign n_28063 = ~x_2415 & ~x_2416;
assign n_28064 = ~x_2417 & ~x_2418;
assign n_28065 =  n_28063 &  n_28064;
assign n_28066 = ~x_2411 & ~x_2412;
assign n_28067 = ~x_2413 & ~x_2414;
assign n_28068 =  n_28066 &  n_28067;
assign n_28069 =  n_28065 &  n_28068;
assign n_28070 = ~x_2423 & ~x_2424;
assign n_28071 = ~x_2425 & ~x_2426;
assign n_28072 =  n_28070 &  n_28071;
assign n_28073 = ~x_2419 & ~x_2420;
assign n_28074 = ~x_2421 & ~x_2422;
assign n_28075 =  n_28073 &  n_28074;
assign n_28076 =  n_28072 &  n_28075;
assign n_28077 =  n_28069 &  n_28076;
assign n_28078 =  n_28062 &  n_28077;
assign n_28079 =  n_28047 &  n_28078;
assign n_28080 =  n_12614 &  n_2303;
assign n_28081 = ~x_2463 & ~x_2464;
assign n_28082 = ~x_2465 & ~x_2466;
assign n_28083 =  n_28081 &  n_28082;
assign n_28084 = ~x_2459 & ~x_2460;
assign n_28085 = ~x_2461 & ~x_2462;
assign n_28086 =  n_28084 &  n_28085;
assign n_28087 =  n_28083 &  n_28086;
assign n_28088 = ~x_2471 & ~x_2472;
assign n_28089 = ~x_2473 & ~x_2474;
assign n_28090 =  n_28088 &  n_28089;
assign n_28091 = ~x_2467 & ~x_2468;
assign n_28092 = ~x_2469 & ~x_2470;
assign n_28093 =  n_28091 &  n_28092;
assign n_28094 =  n_28090 &  n_28093;
assign n_28095 =  n_28087 &  n_28094;
assign n_28096 = ~x_2447 & ~x_2448;
assign n_28097 = ~x_2449 & ~x_2450;
assign n_28098 =  n_28096 &  n_28097;
assign n_28099 = ~x_2443 & ~x_2444;
assign n_28100 = ~x_2445 & ~x_2446;
assign n_28101 =  n_28099 &  n_28100;
assign n_28102 =  n_28098 &  n_28101;
assign n_28103 = ~x_2455 & ~x_2456;
assign n_28104 = ~x_2457 & ~x_2458;
assign n_28105 =  n_28103 &  n_28104;
assign n_28106 = ~x_2451 & ~x_2452;
assign n_28107 = ~x_2453 & ~x_2454;
assign n_28108 =  n_28106 &  n_28107;
assign n_28109 =  n_28105 &  n_28108;
assign n_28110 =  n_28102 &  n_28109;
assign n_28111 =  n_28095 &  n_28110;
assign n_28112 =  n_28080 &  n_28111;
assign n_28113 = ~n_28079 & ~n_28112;
assign n_28114 =  n_4993 &  n_14807;
assign n_28115 =  x_38 &  n_6533;
assign n_28116 =  n_27266 &  n_28115;
assign n_28117 = ~n_28114 & ~n_28116;
assign n_28118 =  n_28113 &  n_28117;
assign n_28119 = ~n_28034 &  n_28035;
assign n_28120 =  n_28118 & ~n_28119;
assign n_28121 =  x_42 &  n_2304;
assign n_28122 =  n_1706 &  n_1180;
assign n_28123 = ~n_28122 & ~n_4639;
assign n_28124 = ~n_13016 &  n_28123;
assign n_28125 = ~n_28121 &  n_28124;
assign n_28126 =  n_2101 &  n_8060;
assign n_28127 = ~n_28034 &  n_28126;
assign n_28128 =  n_28125 & ~n_28127;
assign n_28129 =  n_28120 &  n_28128;
assign n_28130 = ~x_1129 &  n_27810;
assign n_28131 =  n_27973 & ~n_28130;
assign n_28132 =  n_1906 &  n_4056;
assign n_28133 =  n_28131 &  n_28132;
assign n_28134 = ~x_927 & ~x_928;
assign n_28135 = ~x_929 & ~x_930;
assign n_28136 =  n_28134 &  n_28135;
assign n_28137 = ~x_923 & ~x_924;
assign n_28138 = ~x_925 & ~x_926;
assign n_28139 =  n_28137 &  n_28138;
assign n_28140 =  n_28136 &  n_28139;
assign n_28141 = ~x_935 & ~x_936;
assign n_28142 = ~x_937 & ~x_938;
assign n_28143 =  n_28141 &  n_28142;
assign n_28144 = ~x_931 & ~x_932;
assign n_28145 = ~x_933 & ~x_934;
assign n_28146 =  n_28144 &  n_28145;
assign n_28147 =  n_28143 &  n_28146;
assign n_28148 =  n_28140 &  n_28147;
assign n_28149 = ~x_911 & ~x_912;
assign n_28150 = ~x_913 & ~x_914;
assign n_28151 =  n_28149 &  n_28150;
assign n_28152 = ~x_907 & ~x_908;
assign n_28153 = ~x_909 & ~x_910;
assign n_28154 =  n_28152 &  n_28153;
assign n_28155 =  n_28151 &  n_28154;
assign n_28156 = ~x_919 & ~x_920;
assign n_28157 = ~x_921 & ~x_922;
assign n_28158 =  n_28156 &  n_28157;
assign n_28159 = ~x_915 & ~x_916;
assign n_28160 = ~x_917 & ~x_918;
assign n_28161 =  n_28159 &  n_28160;
assign n_28162 =  n_28158 &  n_28161;
assign n_28163 =  n_28155 &  n_28162;
assign n_28164 =  n_28148 &  n_28163;
assign n_28165 =  n_586 &  n_12615;
assign n_28166 = ~n_28164 &  n_28165;
assign n_28167 =  n_186 &  n_6135;
assign n_28168 = ~x_1343 & ~x_1344;
assign n_28169 = ~x_1345 & ~x_1346;
assign n_28170 =  n_28168 &  n_28169;
assign n_28171 = ~x_1339 & ~x_1340;
assign n_28172 = ~x_1341 & ~x_1342;
assign n_28173 =  n_28171 &  n_28172;
assign n_28174 =  n_28170 &  n_28173;
assign n_28175 = ~x_1351 & ~x_1352;
assign n_28176 = ~x_1353 & ~x_1354;
assign n_28177 =  n_28175 &  n_28176;
assign n_28178 = ~x_1347 & ~x_1348;
assign n_28179 = ~x_1349 & ~x_1350;
assign n_28180 =  n_28178 &  n_28179;
assign n_28181 =  n_28177 &  n_28180;
assign n_28182 =  n_28174 &  n_28181;
assign n_28183 = ~x_1327 & ~x_1328;
assign n_28184 = ~x_1329 & ~x_1330;
assign n_28185 =  n_28183 &  n_28184;
assign n_28186 = ~x_1323 & ~x_1324;
assign n_28187 = ~x_1325 & ~x_1326;
assign n_28188 =  n_28186 &  n_28187;
assign n_28189 =  n_28185 &  n_28188;
assign n_28190 = ~x_1335 & ~x_1336;
assign n_28191 = ~x_1337 & ~x_1338;
assign n_28192 =  n_28190 &  n_28191;
assign n_28193 = ~x_1331 & ~x_1332;
assign n_28194 = ~x_1333 & ~x_1334;
assign n_28195 =  n_28193 &  n_28194;
assign n_28196 =  n_28192 &  n_28195;
assign n_28197 =  n_28189 &  n_28196;
assign n_28198 =  n_28182 &  n_28197;
assign n_28199 =  n_28167 &  n_28198;
assign n_28200 = ~n_28166 & ~n_28199;
assign n_28201 =  n_586 &  n_1510;
assign n_28202 =  n_28201 &  n_6330;
assign n_28203 = ~n_22924 & ~n_28202;
assign n_28204 = ~n_7866 & ~n_4994;
assign n_28205 = ~n_7672 &  n_28204;
assign n_28206 =  n_28203 &  n_28205;
assign n_28207 =  n_28200 &  n_28206;
assign n_28208 = ~n_28133 &  n_28207;
assign n_28209 =  n_1 &  n_14808;
assign n_28210 =  n_12614 &  n_12032;
assign n_28211 =  n_3469 &  n_4445;
assign n_28212 = ~n_28210 & ~n_28211;
assign n_28213 = ~n_28209 &  n_28212;
assign n_28214 =  n_10318 &  n_5187;
assign n_28215 = ~n_4252 & ~n_28214;
assign n_28216 =  n_28213 &  n_28215;
assign n_28217 =  n_187 &  n_388;
assign n_28218 =  n_385 &  n_28217;
assign n_28219 =  n_185 &  n_28218;
assign n_28220 = ~n_1317 & ~n_28219;
assign n_28221 = ~n_16721 & ~n_20525;
assign n_28222 =  n_28220 &  n_28221;
assign n_28223 =  n_28216 &  n_28222;
assign n_28224 =  n_28208 &  n_28223;
assign n_28225 =  n_28129 &  n_28224;
assign n_28226 = ~x_1993 &  n_27581;
assign n_28227 = ~x_1994 &  n_28226;
assign n_28228 = ~x_36 &  n_28014;
assign n_28229 = ~n_28227 &  n_28228;
assign n_28230 =  n_23697 &  n_28229;
assign n_28231 = ~x_1130 &  n_28130;
assign n_28232 =  n_27973 & ~n_28231;
assign n_28233 =  x_35 & ~x_36;
assign n_28234 =  n_2100 &  n_8060;
assign n_28235 =  n_28233 &  n_28234;
assign n_28236 =  n_28232 &  n_28235;
assign n_28237 = ~n_28230 & ~n_28236;
assign n_28238 =  n_2499 &  n_24801;
assign n_28239 =  n_28238 &  n_27919;
assign n_28240 =  n_27256 &  n_1313;
assign n_28241 =  n_28240 &  n_1315;
assign n_28242 = ~n_16920 & ~n_28241;
assign n_28243 = ~n_27780 &  n_27835;
assign n_28244 =  n_28242 & ~n_28243;
assign n_28245 =  n_19945 &  n_2296;
assign n_28246 = ~x_1759 & ~x_1760;
assign n_28247 = ~x_1761 & ~x_1762;
assign n_28248 =  n_28246 &  n_28247;
assign n_28249 = ~x_1755 & ~x_1756;
assign n_28250 = ~x_1757 & ~x_1758;
assign n_28251 =  n_28249 &  n_28250;
assign n_28252 =  n_28248 &  n_28251;
assign n_28253 = ~x_1767 & ~x_1768;
assign n_28254 = ~x_1769 & ~x_1770;
assign n_28255 =  n_28253 &  n_28254;
assign n_28256 = ~x_1763 & ~x_1764;
assign n_28257 = ~x_1765 & ~x_1766;
assign n_28258 =  n_28256 &  n_28257;
assign n_28259 =  n_28255 &  n_28258;
assign n_28260 =  n_28252 &  n_28259;
assign n_28261 = ~x_1743 & ~x_1744;
assign n_28262 = ~x_1745 & ~x_1746;
assign n_28263 =  n_28261 &  n_28262;
assign n_28264 = ~x_1739 & ~x_1740;
assign n_28265 = ~x_1741 & ~x_1742;
assign n_28266 =  n_28264 &  n_28265;
assign n_28267 =  n_28263 &  n_28266;
assign n_28268 = ~x_1751 & ~x_1752;
assign n_28269 = ~x_1753 & ~x_1754;
assign n_28270 =  n_28268 &  n_28269;
assign n_28271 = ~x_1747 & ~x_1748;
assign n_28272 = ~x_1749 & ~x_1750;
assign n_28273 =  n_28271 &  n_28272;
assign n_28274 =  n_28270 &  n_28273;
assign n_28275 =  n_28267 &  n_28274;
assign n_28276 =  n_28260 &  n_28275;
assign n_28277 =  n_3 &  n_588;
assign n_28278 = ~n_28276 &  n_28277;
assign n_28279 =  n_6533 &  n_2297;
assign n_28280 = ~x_2399 & ~x_2400;
assign n_28281 = ~x_2401 & ~x_2402;
assign n_28282 =  n_28280 &  n_28281;
assign n_28283 = ~x_2395 & ~x_2396;
assign n_28284 = ~x_2397 & ~x_2398;
assign n_28285 =  n_28283 &  n_28284;
assign n_28286 =  n_28282 &  n_28285;
assign n_28287 = ~x_2407 & ~x_2408;
assign n_28288 = ~x_2409 & ~x_2410;
assign n_28289 =  n_28287 &  n_28288;
assign n_28290 = ~x_2403 & ~x_2404;
assign n_28291 = ~x_2405 & ~x_2406;
assign n_28292 =  n_28290 &  n_28291;
assign n_28293 =  n_28289 &  n_28292;
assign n_28294 =  n_28286 &  n_28293;
assign n_28295 = ~x_2383 & ~x_2384;
assign n_28296 = ~x_2385 & ~x_2386;
assign n_28297 =  n_28295 &  n_28296;
assign n_28298 = ~x_2379 & ~x_2380;
assign n_28299 = ~x_2381 & ~x_2382;
assign n_28300 =  n_28298 &  n_28299;
assign n_28301 =  n_28297 &  n_28300;
assign n_28302 = ~x_2391 & ~x_2392;
assign n_28303 = ~x_2393 & ~x_2394;
assign n_28304 =  n_28302 &  n_28303;
assign n_28305 = ~x_2387 & ~x_2388;
assign n_28306 = ~x_2389 & ~x_2390;
assign n_28307 =  n_28305 &  n_28306;
assign n_28308 =  n_28304 &  n_28307;
assign n_28309 =  n_28301 &  n_28308;
assign n_28310 =  n_28294 &  n_28309;
assign n_28311 =  n_28279 &  n_28310;
assign n_28312 = ~n_28278 & ~n_28311;
assign n_28313 = ~n_28245 &  n_28312;
assign n_28314 =  n_28244 &  n_28313;
assign n_28315 = ~n_28239 &  n_28314;
assign n_28316 =  n_28237 &  n_28315;
assign n_28317 =  n_28225 &  n_28316;
assign n_28318 = ~n_23893 & ~n_16932;
assign n_28319 = ~x_1419 & ~n_27744;
assign n_28320 =  n_586 &  n_3861;
assign n_28321 =  n_6330 &  n_28320;
assign n_28322 = ~n_28319 &  n_28321;
assign n_28323 =  n_28318 & ~n_28322;
assign n_28324 =  n_28164 &  n_28165;
assign n_28325 =  n_1510 &  n_1315;
assign n_28326 =  n_27402 &  n_28325;
assign n_28327 =  n_27266 &  n_28325;
assign n_28328 = ~n_28326 & ~n_28327;
assign n_28329 = ~n_28324 &  n_28328;
assign n_28330 =  n_2 &  n_13006;
assign n_28331 = ~n_28330 & ~n_1513;
assign n_28332 = ~n_21686 &  n_28331;
assign n_28333 =  n_28329 &  n_28332;
assign n_28334 =  n_28323 &  n_28333;
assign n_28335 =  n_587 &  n_3275;
assign n_28336 = ~n_22538 & ~n_28335;
assign n_28337 = ~n_9 &  n_28336;
assign n_28338 =  n_3 &  n_2499;
assign n_28339 = ~n_24220 & ~n_28338;
assign n_28340 =  n_28337 &  n_28339;
assign n_28341 = ~n_27780 &  n_27781;
assign n_28342 = ~n_16925 & ~n_13030;
assign n_28343 = ~n_28341 &  n_28342;
assign n_28344 =  n_28340 &  n_28343;
assign n_28345 =  n_28334 &  n_28344;
assign n_28346 =  n_4993 &  n_2499;
assign n_28347 =  n_388 &  n_28234;
assign n_28348 = ~n_28347 & ~n_6534;
assign n_28349 = ~n_28346 &  n_28348;
assign n_28350 =  n_2 &  n_13015;
assign n_28351 = ~n_15755 & ~n_28350;
assign n_28352 =  n_28349 &  n_28351;
assign n_28353 =  n_783 &  n_1179;
assign n_28354 = ~n_28319 &  n_28353;
assign n_28355 =  n_10520 & ~n_28354;
assign n_28356 =  n_28352 &  n_28355;
assign n_28357 =  n_24801 &  n_27704;
assign n_28358 =  n_3469 &  n_7865;
assign n_28359 = ~x_1311 & ~x_1312;
assign n_28360 = ~x_1313 & ~x_1314;
assign n_28361 =  n_28359 &  n_28360;
assign n_28362 = ~x_1307 & ~x_1308;
assign n_28363 = ~x_1309 & ~x_1310;
assign n_28364 =  n_28362 &  n_28363;
assign n_28365 =  n_28361 &  n_28364;
assign n_28366 = ~x_1319 & ~x_1320;
assign n_28367 = ~x_1321 & ~x_1322;
assign n_28368 =  n_28366 &  n_28367;
assign n_28369 = ~x_1315 & ~x_1316;
assign n_28370 = ~x_1317 & ~x_1318;
assign n_28371 =  n_28369 &  n_28370;
assign n_28372 =  n_28368 &  n_28371;
assign n_28373 =  n_28365 &  n_28372;
assign n_28374 = ~x_1295 & ~x_1296;
assign n_28375 = ~x_1297 & ~x_1298;
assign n_28376 =  n_28374 &  n_28375;
assign n_28377 = ~x_1291 & ~x_1292;
assign n_28378 = ~x_1293 & ~x_1294;
assign n_28379 =  n_28377 &  n_28378;
assign n_28380 =  n_28376 &  n_28379;
assign n_28381 = ~x_1303 & ~x_1304;
assign n_28382 = ~x_1305 & ~x_1306;
assign n_28383 =  n_28381 &  n_28382;
assign n_28384 = ~x_1299 & ~x_1300;
assign n_28385 = ~x_1301 & ~x_1302;
assign n_28386 =  n_28384 &  n_28385;
assign n_28387 =  n_28383 &  n_28386;
assign n_28388 =  n_28380 &  n_28387;
assign n_28389 =  n_28373 &  n_28388;
assign n_28390 =  n_28358 &  n_28389;
assign n_28391 =  n_783 &  n_6135;
assign n_28392 = ~x_1471 & ~x_1472;
assign n_28393 = ~x_1473 & ~x_1474;
assign n_28394 =  n_28392 &  n_28393;
assign n_28395 = ~x_1467 & ~x_1468;
assign n_28396 = ~x_1469 & ~x_1470;
assign n_28397 =  n_28395 &  n_28396;
assign n_28398 =  n_28394 &  n_28397;
assign n_28399 = ~x_1479 & ~x_1480;
assign n_28400 = ~x_1481 & ~x_1482;
assign n_28401 =  n_28399 &  n_28400;
assign n_28402 = ~x_1475 & ~x_1476;
assign n_28403 = ~x_1477 & ~x_1478;
assign n_28404 =  n_28402 &  n_28403;
assign n_28405 =  n_28401 &  n_28404;
assign n_28406 =  n_28398 &  n_28405;
assign n_28407 = ~x_1455 & ~x_1456;
assign n_28408 = ~x_1457 & ~x_1458;
assign n_28409 =  n_28407 &  n_28408;
assign n_28410 = ~x_1451 & ~x_1452;
assign n_28411 = ~x_1453 & ~x_1454;
assign n_28412 =  n_28410 &  n_28411;
assign n_28413 =  n_28409 &  n_28412;
assign n_28414 = ~x_1463 & ~x_1464;
assign n_28415 = ~x_1465 & ~x_1466;
assign n_28416 =  n_28414 &  n_28415;
assign n_28417 = ~x_1459 & ~x_1460;
assign n_28418 = ~x_1461 & ~x_1462;
assign n_28419 =  n_28417 &  n_28418;
assign n_28420 =  n_28416 &  n_28419;
assign n_28421 =  n_28413 &  n_28420;
assign n_28422 =  n_28406 &  n_28421;
assign n_28423 =  n_28391 &  n_28422;
assign n_28424 = ~n_28390 & ~n_28423;
assign n_28425 = ~n_28357 &  n_28424;
assign n_28426 =  x_42 &  n_10521;
assign n_28427 = ~n_28426 & ~n_13869;
assign n_28428 = ~n_22731 & ~n_22072;
assign n_28429 =  n_6533 &  n_3081;
assign n_28430 = ~n_28429 & ~n_1907;
assign n_28431 =  n_28428 &  n_28430;
assign n_28432 =  n_28427 &  n_28431;
assign n_28433 =  n_28425 &  n_28432;
assign n_28434 =  n_28356 &  n_28433;
assign n_28435 =  n_28345 &  n_28434;
assign n_28436 =  n_8254 &  n_1179;
assign n_28437 = ~n_16141 & ~n_28436;
assign n_28438 = ~n_6136 &  n_28437;
assign n_28439 =  n_27256 &  n_27814;
assign n_28440 = ~n_24414 & ~n_28439;
assign n_28441 =  n_1178 &  n_24413;
assign n_28442 = ~n_28441 & ~n_20139;
assign n_28443 =  n_28440 &  n_28442;
assign n_28444 =  n_28438 &  n_28443;
assign n_28445 = ~n_23117 & ~n_21879;
assign n_28446 = ~x_39 &  n_27599;
assign n_28447 =  n_28446 &  n_1315;
assign n_28448 =  n_28445 & ~n_28447;
assign n_28449 =  n_28444 &  n_28448;
assign n_28450 =  n_7 &  n_2302;
assign n_28451 =  n_1 &  n_28450;
assign n_28452 = ~n_28451 & ~n_15948;
assign n_28453 =  n_27413 &  n_1906;
assign n_28454 = ~n_28453 & ~n_13025;
assign n_28455 =  n_28452 &  n_28454;
assign n_28456 = ~n_21493 & ~n_4058;
assign n_28457 =  n_13012 &  n_1510;
assign n_28458 =  n_2296 &  n_28457;
assign n_28459 = ~n_3276 & ~n_28458;
assign n_28460 =  n_28456 &  n_28459;
assign n_28461 =  n_6527 &  n_3;
assign n_28462 = ~n_28461 & ~n_22265;
assign n_28463 =  n_28460 &  n_28462;
assign n_28464 =  n_28455 &  n_28463;
assign n_28465 =  n_28449 &  n_28464;
assign n_28466 =  n_586 & ~n_18429;
assign n_28467 = ~x_42 &  n_23894;
assign n_28468 = ~n_28466 & ~n_28467;
assign n_28469 = ~x_42 &  n_27840;
assign n_28470 =  n_1707 &  n_6527;
assign n_28471 =  n_388 &  n_28022;
assign n_28472 = ~n_28470 & ~n_28471;
assign n_28473 = ~n_28469 &  n_28472;
assign n_28474 =  n_28468 &  n_28473;
assign n_28475 = ~x_2575 & ~x_2576;
assign n_28476 = ~x_2577 & ~x_2578;
assign n_28477 =  n_28475 &  n_28476;
assign n_28478 = ~x_2571 & ~x_2572;
assign n_28479 = ~x_2573 & ~x_2574;
assign n_28480 =  n_28478 &  n_28479;
assign n_28481 =  n_28477 &  n_28480;
assign n_28482 = ~x_2583 & ~x_2584;
assign n_28483 = ~x_2585 & ~x_2586;
assign n_28484 =  n_28482 &  n_28483;
assign n_28485 = ~x_2579 & ~x_2580;
assign n_28486 = ~x_2581 & ~x_2582;
assign n_28487 =  n_28485 &  n_28486;
assign n_28488 =  n_28484 &  n_28487;
assign n_28489 =  n_28481 &  n_28488;
assign n_28490 =  n_3469 &  n_28489;
assign n_28491 = ~x_2591 & ~x_2592;
assign n_28492 = ~x_2593 & ~x_2594;
assign n_28493 =  n_28491 &  n_28492;
assign n_28494 = ~x_2587 & ~x_2588;
assign n_28495 = ~x_2589 & ~x_2590;
assign n_28496 =  n_28494 &  n_28495;
assign n_28497 =  n_28493 &  n_28496;
assign n_28498 = ~x_2599 & ~x_2600;
assign n_28499 = ~x_2601 & ~x_2602;
assign n_28500 =  n_28498 &  n_28499;
assign n_28501 = ~x_2595 & ~x_2596;
assign n_28502 = ~x_2597 & ~x_2598;
assign n_28503 =  n_28501 &  n_28502;
assign n_28504 =  n_28500 &  n_28503;
assign n_28505 =  n_28497 &  n_28504;
assign n_28506 =  n_23891 &  n_28505;
assign n_28507 =  n_28490 &  n_28506;
assign n_28508 =  n_1906 &  n_27403;
assign n_28509 = ~n_28507 & ~n_28508;
assign n_28510 = ~n_20332 & ~n_13021;
assign n_28511 =  n_10318 &  n_13006;
assign n_28512 =  n_8818 &  n_983;
assign n_28513 = ~n_28511 & ~n_28512;
assign n_28514 =  n_28510 &  n_28513;
assign n_28515 =  n_28509 &  n_28514;
assign n_28516 =  n_28474 &  n_28515;
assign n_28517 =  n_28465 &  n_28516;
assign n_28518 =  n_12420 &  n_27971;
assign n_28519 =  n_3664 &  n_4;
assign n_28520 =  n_28011 &  n_28519;
assign n_28521 = ~n_28518 & ~n_28520;
assign n_28522 = ~x_38 &  n_27274;
assign n_28523 =  n_8254 &  n_28522;
assign n_28524 =  n_1314 &  n_5191;
assign n_28525 =  n_28201 &  n_27274;
assign n_28526 = ~n_28524 & ~n_28525;
assign n_28527 = ~n_28523 &  n_28526;
assign n_28528 =  x_38 &  n_27258;
assign n_28529 =  n_1707 &  n_28528;
assign n_28530 = ~n_28529 & ~n_24995;
assign n_28531 =  n_28527 &  n_28530;
assign n_28532 =  n_28521 &  n_28531;
assign n_28533 =  n_585 &  n_13006;
assign n_28534 = ~n_28533 & ~n_24607;
assign n_28535 =  n_27257 &  n_187;
assign n_28536 =  n_28535 &  n_1906;
assign n_28537 =  n_24801 &  n_3275;
assign n_28538 =  n_10318 &  n_10518;
assign n_28539 = ~n_28537 & ~n_28538;
assign n_28540 = ~n_28536 &  n_28539;
assign n_28541 =  n_28534 &  n_28540;
assign n_28542 = ~n_18440 & ~n_24802;
assign n_28543 =  n_1315 &  n_13006;
assign n_28544 = ~n_13013 & ~n_28543;
assign n_28545 =  n_28542 &  n_28544;
assign n_28546 =  n_28541 &  n_28545;
assign n_28547 =  n_4992 &  n_28218;
assign n_28548 = ~n_2693 & ~n_28547;
assign n_28549 =  n_3664 &  n_14807;
assign n_28550 =  n_10318 &  n_8802;
assign n_28551 =  n_4992 &  n_13020;
assign n_28552 = ~n_28550 & ~n_28551;
assign n_28553 = ~n_28549 &  n_28552;
assign n_28554 =  n_28548 &  n_28553;
assign n_28555 =  n_28546 &  n_28554;
assign n_28556 =  n_28532 &  n_28555;
assign n_28557 =  n_28517 &  n_28556;
assign n_28558 =  n_28435 &  n_28557;
assign n_28559 =  n_28317 &  n_28558;
assign n_28560 =  n_28046 &  n_28559;
assign n_28561 =  n_27939 &  n_28560;
assign n_28562 = ~n_27553 &  n_28561;
assign n_28563 = ~n_27426 &  n_28562;
assign n_28564 =  n_27254 &  n_27417;
assign n_28565 =  n_2886 &  n_27402;
assign n_28566 =  n_10318 &  n_28565;
assign n_28567 =  n_27254 &  n_28566;
assign n_28568 = ~n_28564 & ~n_28567;
assign n_28569 =  n_28563 &  n_28568;
assign n_28570 =  n_8818 &  n_27260;
assign n_28571 = ~n_27254 &  n_27404;
assign n_28572 = ~n_27254 &  n_27414;
assign n_28573 = ~n_28571 & ~n_28572;
assign n_28574 = ~n_28570 &  n_28573;
assign n_28575 =  n_28569 &  n_28574;
assign n_28576 =  n_27421 &  n_28575;
assign n_28577 =  n_27272 &  n_28576;
assign n_28578 =  n_27266 &  n_25774;
assign n_28579 = ~n_27399 &  n_28578;
assign n_28580 =  n_4992 &  n_28240;
assign n_28581 = ~n_27399 &  n_28580;
assign n_28582 = ~x_40 &  n_28581;
assign n_28583 = ~n_28579 & ~n_28582;
assign n_28584 =  n_8060 &  n_27411;
assign n_28585 =  x_38 &  n_27402;
assign n_28586 =  n_8818 &  n_28585;
assign n_28587 =  n_27254 &  n_28586;
assign n_28588 = ~n_28584 & ~n_28587;
assign n_28589 =  n_12420 &  n_28535;
assign n_28590 = ~n_27399 &  n_28589;
assign n_28591 =  x_40 &  n_28581;
assign n_28592 = ~n_28590 & ~n_28591;
assign n_28593 =  n_28588 &  n_28592;
assign n_28594 =  n_28583 &  n_28593;
assign n_28595 =  n_27254 &  n_27599;
assign n_28596 =  n_8818 &  n_28595;
assign n_28597 =  n_28595 &  n_3664;
assign n_28598 = ~n_28596 & ~n_28597;
assign n_28599 =  n_27262 &  n_2;
assign n_28600 =  n_4993 &  n_27424;
assign n_28601 = ~n_28599 & ~n_28600;
assign n_28602 =  n_3 &  n_28522;
assign n_28603 =  n_28601 & ~n_28602;
assign n_28604 = ~n_27399 & ~n_28603;
assign n_28605 =  n_3664 &  n_27406;
assign n_28606 =  n_27254 &  n_28605;
assign n_28607 = ~n_28446 & ~n_27593;
assign n_28608 =  n_4992 & ~n_28607;
assign n_28609 = ~n_27399 &  n_28608;
assign n_28610 = ~n_28606 & ~n_28609;
assign n_28611 = ~n_28604 &  n_28610;
assign n_28612 =  n_28598 &  n_28611;
assign n_28613 = ~n_27254 &  n_27267;
assign n_28614 =  n_3664 &  n_28613;
assign n_28615 =  n_8818 &  n_28613;
assign n_28616 = ~n_28614 & ~n_28615;
assign n_28617 =  n_586 &  n_27263;
assign n_28618 =  n_27400 &  n_27402;
assign n_28619 = ~n_28617 & ~n_28618;
assign n_28620 =  n_28616 &  n_28619;
assign n_28621 =  n_28612 &  n_28620;
assign n_28622 =  n_28594 &  n_28621;
assign n_28623 =  n_28577 &  n_28622;
assign n_28624 = ~n_27129 &  n_28623;
assign n_28625 = ~n_26679 &  n_28624;
assign n_28626 =  n_26228 &  n_28625;
assign n_28627 =  x_42 &  n_28626;
assign n_28628 = ~x_42 & ~n_28626;
assign n_28629 = ~n_28627 & ~n_28628;
assign n_28630 =  n_26229 & ~n_26678;
assign n_28631 = ~n_27129 &  n_28592;
assign n_28632 = ~n_27254 &  n_27425;
assign n_28633 = ~n_28614 & ~n_28632;
assign n_28634 = ~n_27254 &  n_27259;
assign n_28635 =  n_3664 &  n_28634;
assign n_28636 =  n_13012 &  n_27411;
assign n_28637 = ~n_28635 & ~n_28636;
assign n_28638 =  n_28633 &  n_28637;
assign n_28639 =  n_28537 & ~n_28029;
assign n_28640 =  n_28538 & ~n_27703;
assign n_28641 = ~n_27826 & ~n_28640;
assign n_28642 = ~n_28639 &  n_28641;
assign n_28643 = ~n_28036 &  n_28642;
assign n_28644 =  n_6533 &  n_4445;
assign n_28645 = ~n_28357 & ~n_28644;
assign n_28646 =  n_28645 & ~n_28551;
assign n_28647 =  n_27422 &  n_28201;
assign n_28648 =  n_28017 &  n_28647;
assign n_28649 = ~n_28648 & ~n_27972;
assign n_28650 =  n_28646 &  n_28649;
assign n_28651 =  n_27935 &  n_28650;
assign n_28652 =  n_28643 &  n_28651;
assign n_28653 =  n_24413 &  n_28023;
assign n_28654 = ~x_543 & ~x_544;
assign n_28655 = ~x_545 & ~x_546;
assign n_28656 =  n_28654 &  n_28655;
assign n_28657 = ~x_539 & ~x_540;
assign n_28658 = ~x_541 & ~x_542;
assign n_28659 =  n_28657 &  n_28658;
assign n_28660 =  n_28656 &  n_28659;
assign n_28661 = ~x_551 & ~x_552;
assign n_28662 = ~x_553 & ~x_554;
assign n_28663 =  n_28661 &  n_28662;
assign n_28664 = ~x_547 & ~x_548;
assign n_28665 = ~x_549 & ~x_550;
assign n_28666 =  n_28664 &  n_28665;
assign n_28667 =  n_28663 &  n_28666;
assign n_28668 =  n_28660 &  n_28667;
assign n_28669 = ~x_527 & ~x_528;
assign n_28670 = ~x_529 & ~x_530;
assign n_28671 =  n_28669 &  n_28670;
assign n_28672 = ~x_523 & ~x_524;
assign n_28673 = ~x_525 & ~x_526;
assign n_28674 =  n_28672 &  n_28673;
assign n_28675 =  n_28671 &  n_28674;
assign n_28676 = ~x_535 & ~x_536;
assign n_28677 = ~x_537 & ~x_538;
assign n_28678 =  n_28676 &  n_28677;
assign n_28679 = ~x_531 & ~x_532;
assign n_28680 = ~x_533 & ~x_534;
assign n_28681 =  n_28679 &  n_28680;
assign n_28682 =  n_28678 &  n_28681;
assign n_28683 =  n_28675 &  n_28682;
assign n_28684 =  n_28668 &  n_28683;
assign n_28685 =  n_1707 &  n_2499;
assign n_28686 =  n_28684 &  n_28685;
assign n_28687 = ~n_28653 & ~n_28686;
assign n_28688 = ~n_28684 &  n_28685;
assign n_28689 = ~n_27834 & ~n_28688;
assign n_28690 =  n_28687 &  n_28689;
assign n_28691 =  n_28652 &  n_28690;
assign n_28692 =  n_10318 &  n_3862;
assign n_28693 = ~n_14817 & ~n_28692;
assign n_28694 =  n_6533 &  n_28217;
assign n_28695 = ~n_28694 & ~n_18440;
assign n_28696 =  n_28693 &  n_28695;
assign n_28697 =  n_3081 &  n_24801;
assign n_28698 = ~n_25775 & ~n_8256;
assign n_28699 = ~n_28697 &  n_28698;
assign n_28700 =  n_14807 &  n_980;
assign n_28701 =  n_3664 &  n_390;
assign n_28702 = ~n_28700 & ~n_28701;
assign n_28703 =  n_28699 &  n_28702;
assign n_28704 =  n_28696 &  n_28703;
assign n_28705 = ~n_16919 & ~n_8813;
assign n_28706 =  n_1315 &  n_8803;
assign n_28707 = ~n_10516 & ~n_28706;
assign n_28708 =  n_28705 &  n_28707;
assign n_28709 = ~n_27916 & ~n_27835;
assign n_28710 = ~n_28338 & ~n_27588;
assign n_28711 =  n_28709 &  n_28710;
assign n_28712 =  n_28708 &  n_28711;
assign n_28713 =  n_28704 &  n_28712;
assign n_28714 = ~n_28447 & ~n_28507;
assign n_28715 =  n_979 &  n_28218;
assign n_28716 =  n_6533 &  n_8;
assign n_28717 =  n_14807 &  n_1707;
assign n_28718 = ~n_28716 & ~n_28717;
assign n_28719 = ~n_28715 &  n_28718;
assign n_28720 =  n_28714 &  n_28719;
assign n_28721 = ~n_7479 & ~n_589;
assign n_28722 =  n_6533 &  n_4057;
assign n_28723 =  n_1511 &  n_28325;
assign n_28724 = ~n_28722 & ~n_28723;
assign n_28725 = ~n_8819 &  n_28724;
assign n_28726 =  n_28721 &  n_28725;
assign n_28727 =  n_27424 &  n_1906;
assign n_28728 =  n_1709 &  n_24801;
assign n_28729 = ~n_28727 & ~n_28728;
assign n_28730 = ~n_28327 & ~n_14812;
assign n_28731 =  n_28729 &  n_28730;
assign n_28732 =  n_28726 &  n_28731;
assign n_28733 =  n_28720 &  n_28732;
assign n_28734 =  n_28713 &  n_28733;
assign n_28735 = ~n_27598 & ~n_2888;
assign n_28736 =  n_28047 & ~n_28078;
assign n_28737 = ~n_28736 & ~n_27876;
assign n_28738 =  n_28735 &  n_28737;
assign n_28739 =  n_27423 &  n_28325;
assign n_28740 = ~n_28739 & ~n_27912;
assign n_28741 =  n_12614 &  n_23892;
assign n_28742 =  n_27811 &  n_28741;
assign n_28743 =  n_28740 & ~n_28742;
assign n_28744 =  n_28738 &  n_28743;
assign n_28745 = ~n_28038 & ~n_25320;
assign n_28746 =  n_28745 & ~n_13016;
assign n_28747 =  n_3663 &  n_6527;
assign n_28748 = ~n_10522 & ~n_28747;
assign n_28749 =  n_28746 &  n_28748;
assign n_28750 =  n_1707 &  n_2101;
assign n_28751 = ~n_20139 & ~n_28750;
assign n_28752 = ~x_41 &  n_13020;
assign n_28753 =  n_28751 & ~n_28752;
assign n_28754 =  n_1706 &  n_12615;
assign n_28755 = ~n_28754 &  n_27707;
assign n_28756 =  n_28753 &  n_28755;
assign n_28757 =  n_28749 &  n_28756;
assign n_28758 =  x_37 &  n_7;
assign n_28759 =  n_6530 &  n_28758;
assign n_28760 =  n_14807 &  n_6533;
assign n_28761 = ~n_6137 & ~n_28760;
assign n_28762 = ~n_28759 &  n_28761;
assign n_28763 =  n_28113 &  n_28762;
assign n_28764 =  n_28757 &  n_28763;
assign n_28765 =  n_28744 &  n_28764;
assign n_28766 =  n_28734 &  n_28765;
assign n_28767 =  x_42 &  n_2300;
assign n_28768 = ~n_28458 & ~n_28767;
assign n_28769 =  n_28768 & ~n_3665;
assign n_28770 =  n_1707 &  n_8;
assign n_28771 =  n_6533 &  n_28522;
assign n_28772 = ~n_28770 & ~n_28771;
assign n_28773 =  n_8254 &  n_27416;
assign n_28774 =  n_586 &  n_14808;
assign n_28775 = ~n_28773 & ~n_28774;
assign n_28776 =  n_28772 &  n_28775;
assign n_28777 =  n_28769 &  n_28776;
assign n_28778 =  n_27258 &  n_28325;
assign n_28779 = ~n_28778 & ~n_28467;
assign n_28780 =  n_27258 &  n_6533;
assign n_28781 =  x_38 &  n_28780;
assign n_28782 =  n_1906 &  n_28522;
assign n_28783 = ~n_28781 & ~n_28782;
assign n_28784 =  n_28779 &  n_28783;
assign n_28785 = ~n_16141 &  n_28332;
assign n_28786 =  n_28784 &  n_28785;
assign n_28787 =  n_28777 &  n_28786;
assign n_28788 =  n_1708 &  n_27820;
assign n_28789 = ~n_28788 & ~n_15948;
assign n_28790 = ~x_2175 & ~x_2176;
assign n_28791 = ~x_2177 & ~x_2178;
assign n_28792 =  n_28790 &  n_28791;
assign n_28793 = ~x_2171 & ~x_2172;
assign n_28794 = ~x_2173 & ~x_2174;
assign n_28795 =  n_28793 &  n_28794;
assign n_28796 =  n_28792 &  n_28795;
assign n_28797 = ~x_2183 & ~x_2184;
assign n_28798 = ~x_2185 & ~x_2186;
assign n_28799 =  n_28797 &  n_28798;
assign n_28800 = ~x_2179 & ~x_2180;
assign n_28801 = ~x_2181 & ~x_2182;
assign n_28802 =  n_28800 &  n_28801;
assign n_28803 =  n_28799 &  n_28802;
assign n_28804 =  n_28796 &  n_28803;
assign n_28805 = ~x_2159 & ~x_2160;
assign n_28806 = ~x_2161 & ~x_2162;
assign n_28807 =  n_28805 &  n_28806;
assign n_28808 = ~x_2155 & ~x_2156;
assign n_28809 = ~x_2157 & ~x_2158;
assign n_28810 =  n_28808 &  n_28809;
assign n_28811 =  n_28807 &  n_28810;
assign n_28812 = ~x_2167 & ~x_2168;
assign n_28813 = ~x_2169 & ~x_2170;
assign n_28814 =  n_28812 &  n_28813;
assign n_28815 = ~x_2163 & ~x_2164;
assign n_28816 = ~x_2165 & ~x_2166;
assign n_28817 =  n_28815 &  n_28816;
assign n_28818 =  n_28814 &  n_28817;
assign n_28819 =  n_28811 &  n_28818;
assign n_28820 =  n_28804 &  n_28819;
assign n_28821 =  n_28436 & ~n_28820;
assign n_28822 =  n_28789 & ~n_28821;
assign n_28823 =  n_2 &  n_14808;
assign n_28824 =  n_1315 &  n_6332;
assign n_28825 = ~n_28543 & ~n_28824;
assign n_28826 = ~n_28823 &  n_28825;
assign n_28827 =  n_28822 &  n_28826;
assign n_28828 =  n_1315 &  n_4251;
assign n_28829 =  n_6330 &  n_784;
assign n_28830 = ~n_28828 & ~n_28829;
assign n_28831 = ~n_27839 &  n_28830;
assign n_28832 = ~x_41 &  n_13868;
assign n_28833 = ~n_8818 & ~n_1707;
assign n_28834 =  n_191 & ~n_28833;
assign n_28835 = ~n_28834 & ~n_8824;
assign n_28836 = ~n_28832 &  n_28835;
assign n_28837 =  n_28831 &  n_28836;
assign n_28838 =  n_28827 &  n_28837;
assign n_28839 = ~x_42 &  n_28533;
assign n_28840 = ~n_28121 &  n_28205;
assign n_28841 = ~n_28839 &  n_28840;
assign n_28842 = ~n_28133 &  n_28841;
assign n_28843 =  n_28838 &  n_28842;
assign n_28844 =  n_28787 &  n_28843;
assign n_28845 =  n_28766 &  n_28844;
assign n_28846 =  n_8255 &  n_28229;
assign n_28847 =  n_1706 &  n_27585;
assign n_28848 = ~n_27925 & ~n_28847;
assign n_28849 =  n_1707 &  n_12226;
assign n_28850 =  n_28510 & ~n_28849;
assign n_28851 =  n_28848 &  n_28850;
assign n_28852 = ~n_27587 &  n_28851;
assign n_28853 = ~n_28846 &  n_28852;
assign n_28854 = ~n_13030 & ~n_28469;
assign n_28855 =  x_42 &  n_24607;
assign n_28856 = ~n_28855 & ~n_13025;
assign n_28857 =  n_28854 &  n_28856;
assign n_28858 = ~n_28119 &  n_28857;
assign n_28859 =  n_27273 &  n_8255;
assign n_28860 = ~n_27978 & ~n_28859;
assign n_28861 =  n_28858 &  n_28860;
assign n_28862 =  n_28853 &  n_28861;
assign n_28863 =  n_27267 &  n_8254;
assign n_28864 = ~n_28863 & ~n_27602;
assign n_28865 =  n_28080 & ~n_28111;
assign n_28866 =  n_28358 & ~n_28389;
assign n_28867 = ~n_28865 & ~n_28866;
assign n_28868 =  n_28864 &  n_28867;
assign n_28869 =  n_28868 &  n_28352;
assign n_28870 = ~n_28536 & ~n_23310;
assign n_28871 = ~n_16927 &  n_28870;
assign n_28872 = ~x_42 &  n_23893;
assign n_28873 =  n_28871 & ~n_28872;
assign n_28874 = ~n_9 & ~n_392;
assign n_28875 = ~n_13013 & ~n_16925;
assign n_28876 =  n_28874 &  n_28875;
assign n_28877 =  n_28873 &  n_28876;
assign n_28878 =  n_28869 &  n_28877;
assign n_28879 = ~x_1407 & ~x_1408;
assign n_28880 = ~x_1409 & ~x_1410;
assign n_28881 =  n_28879 &  n_28880;
assign n_28882 = ~x_1403 & ~x_1404;
assign n_28883 = ~x_1405 & ~x_1406;
assign n_28884 =  n_28882 &  n_28883;
assign n_28885 =  n_28881 &  n_28884;
assign n_28886 = ~x_1415 & ~x_1416;
assign n_28887 = ~x_1417 & ~x_1418;
assign n_28888 =  n_28886 &  n_28887;
assign n_28889 = ~x_1411 & ~x_1412;
assign n_28890 = ~x_1413 & ~x_1414;
assign n_28891 =  n_28889 &  n_28890;
assign n_28892 =  n_28888 &  n_28891;
assign n_28893 =  n_28885 &  n_28892;
assign n_28894 = ~x_1391 & ~x_1392;
assign n_28895 = ~x_1393 & ~x_1394;
assign n_28896 =  n_28894 &  n_28895;
assign n_28897 = ~x_1387 & ~x_1388;
assign n_28898 = ~x_1389 & ~x_1390;
assign n_28899 =  n_28897 &  n_28898;
assign n_28900 =  n_28896 &  n_28899;
assign n_28901 = ~x_1399 & ~x_1400;
assign n_28902 = ~x_1401 & ~x_1402;
assign n_28903 =  n_28901 &  n_28902;
assign n_28904 = ~x_1395 & ~x_1396;
assign n_28905 = ~x_1397 & ~x_1398;
assign n_28906 =  n_28904 &  n_28905;
assign n_28907 =  n_28903 &  n_28906;
assign n_28908 =  n_28900 &  n_28907;
assign n_28909 =  n_28893 &  n_28908;
assign n_28910 =  n_6532 &  n_28909;
assign n_28911 =  n_8254 &  n_28910;
assign n_28912 =  n_12420 &  n_28910;
assign n_28913 =  n_10318 &  n_10320;
assign n_28914 =  n_783 &  n_1709;
assign n_28915 =  n_1906 &  n_28217;
assign n_28916 = ~n_28914 & ~n_28915;
assign n_28917 = ~n_28913 &  n_28916;
assign n_28918 = ~n_28912 &  n_28917;
assign n_28919 = ~n_28911 &  n_28918;
assign n_28920 =  n_28919 & ~n_28230;
assign n_28921 =  n_28878 &  n_28920;
assign n_28922 =  n_28862 &  n_28921;
assign n_28923 =  n_28845 &  n_28922;
assign n_28924 =  n_27820 &  n_27747;
assign n_28925 = ~n_28924 & ~n_27749;
assign n_28926 =  n_27748 &  n_27821;
assign n_28927 =  n_6533 &  n_2499;
assign n_28928 =  n_28927 &  n_28684;
assign n_28929 = ~n_28926 & ~n_28928;
assign n_28930 =  n_28927 & ~n_28684;
assign n_28931 = ~n_28930 & ~n_28341;
assign n_28932 =  n_28931 &  n_27818;
assign n_28933 =  n_28929 &  n_28932;
assign n_28934 =  n_28925 &  n_28933;
assign n_28935 = ~n_28226 &  n_28014;
assign n_28936 =  n_27422 &  n_28320;
assign n_28937 =  n_28935 &  n_28936;
assign n_28938 = ~n_28518 & ~n_28937;
assign n_28939 =  n_1311 &  n_28320;
assign n_28940 =  n_28935 &  n_28939;
assign n_28941 =  n_28938 & ~n_28940;
assign n_28942 =  n_28022 &  n_27833;
assign n_28943 =  n_1707 &  n_27403;
assign n_28944 =  n_12420 &  n_23891;
assign n_28945 = ~n_24220 & ~n_28944;
assign n_28946 = ~n_28943 &  n_28945;
assign n_28947 =  n_28279 & ~n_28310;
assign n_28948 =  n_1315 &  n_28450;
assign n_28949 =  n_27256 &  n_1315;
assign n_28950 =  n_27813 &  n_28949;
assign n_28951 = ~n_28948 & ~n_28950;
assign n_28952 = ~n_28529 &  n_28951;
assign n_28953 = ~n_28947 &  n_28952;
assign n_28954 =  n_28946 &  n_28953;
assign n_28955 =  n_28238 & ~n_27919;
assign n_28956 = ~n_28955 &  n_28313;
assign n_28957 =  n_28954 &  n_28956;
assign n_28958 = ~n_28942 &  n_28957;
assign n_28959 =  n_28941 &  n_28958;
assign n_28960 =  n_28934 &  n_28959;
assign n_28961 =  n_28923 &  n_28960;
assign n_28962 =  n_28691 &  n_28961;
assign n_28963 = ~n_27408 &  n_28962;
assign n_28964 = ~n_28609 & ~n_28604;
assign n_28965 =  n_28963 &  n_28964;
assign n_28966 = ~n_27401 & ~n_28618;
assign n_28967 =  n_28965 &  n_28966;
assign n_28968 =  n_28583 &  n_28967;
assign n_28969 =  n_28638 &  n_28968;
assign n_28970 =  n_28631 &  n_28969;
assign n_28971 = ~n_28630 &  n_28970;
assign n_28972 =  x_41 & ~n_28971;
assign n_28973 = ~x_41 &  n_28971;
assign n_28974 = ~n_28972 & ~n_28973;
assign n_28975 = ~n_27639 & ~n_28036;
assign n_28976 =  n_28975 &  n_27921;
assign n_28977 =  n_27929 &  n_28976;
assign n_28978 = ~n_18440 & ~n_1710;
assign n_28979 = ~n_16927 &  n_28978;
assign n_28980 = ~n_4252 & ~n_20525;
assign n_28981 =  n_28980 & ~n_28466;
assign n_28982 =  n_28979 &  n_28981;
assign n_28983 = ~n_28821 & ~n_13474;
assign n_28984 =  n_28983 &  n_28867;
assign n_28985 =  n_28982 &  n_28984;
assign n_28986 =  n_3469 &  n_28522;
assign n_28987 =  n_2 &  n_5187;
assign n_28988 = ~n_28986 & ~n_28987;
assign n_28989 =  n_7 &  n_8255;
assign n_28990 =  n_28730 & ~n_28989;
assign n_28991 =  n_28988 &  n_28990;
assign n_28992 =  n_28113 &  n_28768;
assign n_28993 =  n_28991 &  n_28992;
assign n_28994 =  n_28985 &  n_28993;
assign n_28995 = ~n_28133 & ~n_27817;
assign n_28996 = ~n_28230 &  n_28995;
assign n_28997 =  n_28994 &  n_28996;
assign n_28998 =  n_28977 &  n_28997;
assign n_28999 =  n_1904 &  n_186;
assign n_29000 = ~n_28999 & ~n_28742;
assign n_29001 =  n_28031 &  n_29000;
assign n_29002 =  n_29001 &  n_28689;
assign n_29003 =  n_28998 &  n_29002;
assign n_29004 = ~n_28942 &  n_28925;
assign n_29005 = ~n_27978 & ~n_28739;
assign n_29006 =  n_28649 &  n_29005;
assign n_29007 =  n_29006 &  n_28941;
assign n_29008 =  n_29004 &  n_29007;
assign n_29009 =  n_27877 &  n_27908;
assign n_29010 = ~n_29009 & ~n_28439;
assign n_29011 = ~n_28782 &  n_29010;
assign n_29012 = ~n_27671 &  n_29011;
assign n_29013 = ~n_12227 & ~n_13025;
assign n_29014 =  n_3858 &  n_12032;
assign n_29015 = ~n_13021 & ~n_29014;
assign n_29016 =  n_29013 &  n_29015;
assign n_29017 =  n_29016 &  n_28125;
assign n_29018 =  n_29012 &  n_29017;
assign n_29019 = ~n_28322 & ~n_28533;
assign n_29020 =  n_28931 &  n_29019;
assign n_29021 =  n_8254 &  n_28528;
assign n_29022 =  n_190 &  n_28320;
assign n_29023 = ~n_29021 & ~n_29022;
assign n_29024 = ~x_1727 & ~x_1728;
assign n_29025 = ~x_1729 & ~x_1730;
assign n_29026 =  n_29024 &  n_29025;
assign n_29027 = ~x_1723 & ~x_1724;
assign n_29028 = ~x_1725 & ~x_1726;
assign n_29029 =  n_29027 &  n_29028;
assign n_29030 =  n_29026 &  n_29029;
assign n_29031 = ~x_1735 & ~x_1736;
assign n_29032 = ~x_1737 & ~x_1738;
assign n_29033 =  n_29031 &  n_29032;
assign n_29034 = ~x_1731 & ~x_1732;
assign n_29035 = ~x_1733 & ~x_1734;
assign n_29036 =  n_29034 &  n_29035;
assign n_29037 =  n_29033 &  n_29036;
assign n_29038 =  n_29030 &  n_29037;
assign n_29039 = ~x_1711 & ~x_1712;
assign n_29040 = ~x_1713 & ~x_1714;
assign n_29041 =  n_29039 &  n_29040;
assign n_29042 = ~x_1707 & ~x_1708;
assign n_29043 = ~x_1709 & ~x_1710;
assign n_29044 =  n_29042 &  n_29043;
assign n_29045 =  n_29041 &  n_29044;
assign n_29046 = ~x_1719 & ~x_1720;
assign n_29047 = ~x_1721 & ~x_1722;
assign n_29048 =  n_29046 &  n_29047;
assign n_29049 = ~x_1715 & ~x_1716;
assign n_29050 = ~x_1717 & ~x_1718;
assign n_29051 =  n_29049 &  n_29050;
assign n_29052 =  n_29048 &  n_29051;
assign n_29053 =  n_29045 &  n_29052;
assign n_29054 =  n_29038 &  n_29053;
assign n_29055 =  n_28915 & ~n_29054;
assign n_29056 = ~n_29055 & ~n_27711;
assign n_29057 =  n_29023 &  n_29056;
assign n_29058 = ~n_3470 & ~n_589;
assign n_29059 = ~n_3082 &  n_29058;
assign n_29060 =  n_27910 &  n_29059;
assign n_29061 =  n_29057 &  n_29060;
assign n_29062 =  n_29020 &  n_29061;
assign n_29063 =  n_29018 &  n_29062;
assign n_29064 =  n_6 &  n_27814;
assign n_29065 = ~n_29064 & ~n_28846;
assign n_29066 = ~n_28127 & ~n_28955;
assign n_29067 =  n_28244 &  n_29066;
assign n_29068 =  n_29065 &  n_29067;
assign n_29069 =  n_29063 &  n_29068;
assign n_29070 =  n_27259 &  n_8254;
assign n_29071 = ~n_29070 & ~n_28219;
assign n_29072 =  n_6330 &  n_6530;
assign n_29073 = ~n_27588 & ~n_29072;
assign n_29074 =  n_186 &  n_983;
assign n_29075 = ~n_28543 & ~n_29074;
assign n_29076 =  n_29073 &  n_29075;
assign n_29077 =  n_29071 &  n_29076;
assign n_29078 =  n_186 &  n_28585;
assign n_29079 = ~n_29078 & ~n_28774;
assign n_29080 =  n_186 &  n_27416;
assign n_29081 = ~n_29080 & ~n_28586;
assign n_29082 =  n_29079 &  n_29081;
assign n_29083 =  n_29077 &  n_29082;
assign n_29084 = ~x_42 &  n_28451;
assign n_29085 = ~n_29084 & ~n_28311;
assign n_29086 = ~n_28913 & ~n_28727;
assign n_29087 =  n_29086 & ~n_28166;
assign n_29088 =  n_29085 &  n_29087;
assign n_29089 =  n_27424 &  n_8254;
assign n_29090 = ~n_29089 & ~n_8813;
assign n_29091 = ~n_15755 &  n_29090;
assign n_29092 =  n_6533 &  n_28585;
assign n_29093 = ~n_10517 & ~n_29092;
assign n_29094 =  n_29091 &  n_29093;
assign n_29095 =  n_29088 &  n_29094;
assign n_29096 =  n_29083 &  n_29095;
assign n_29097 =  n_3469 &  n_14807;
assign n_29098 = ~n_16932 & ~n_29097;
assign n_29099 = ~n_12809 & ~n_12616;
assign n_29100 =  n_29098 &  n_29099;
assign n_29101 =  n_980 &  n_390;
assign n_29102 = ~n_29101 & ~n_28347;
assign n_29103 = ~n_5197 & ~n_28780;
assign n_29104 =  n_29102 &  n_29103;
assign n_29105 =  n_29100 &  n_29104;
assign n_29106 = ~n_1181 & ~n_24027;
assign n_29107 = ~n_2500 &  n_29106;
assign n_29108 = ~n_28912 &  n_29107;
assign n_29109 =  n_29105 &  n_29108;
assign n_29110 = ~n_21493 & ~n_28202;
assign n_29111 = ~n_27267 & ~n_27424;
assign n_29112 =  n_186 & ~n_29111;
assign n_29113 =  n_29110 & ~n_29112;
assign n_29114 = ~n_28700 & ~n_28470;
assign n_29115 = ~n_28461 & ~n_28429;
assign n_29116 =  n_29114 &  n_29115;
assign n_29117 =  n_29113 &  n_29116;
assign n_29118 = ~n_28788 & ~n_2888;
assign n_29119 = ~n_22731 &  n_29118;
assign n_29120 = ~n_23503 & ~n_28210;
assign n_29121 =  n_29119 &  n_29120;
assign n_29122 =  n_1707 &  n_28522;
assign n_29123 = ~n_13667 & ~n_8824;
assign n_29124 = ~n_6136 &  n_29123;
assign n_29125 = ~n_29122 &  n_29124;
assign n_29126 =  n_29121 &  n_29125;
assign n_29127 =  n_29117 &  n_29126;
assign n_29128 =  n_29109 &  n_29127;
assign n_29129 =  n_29096 &  n_29128;
assign n_29130 = ~x_1375 & ~x_1376;
assign n_29131 = ~x_1377 & ~x_1378;
assign n_29132 =  n_29130 &  n_29131;
assign n_29133 = ~x_1371 & ~x_1372;
assign n_29134 = ~x_1373 & ~x_1374;
assign n_29135 =  n_29133 &  n_29134;
assign n_29136 =  n_29132 &  n_29135;
assign n_29137 = ~x_1383 & ~x_1384;
assign n_29138 = ~x_1385 & ~x_1386;
assign n_29139 =  n_29137 &  n_29138;
assign n_29140 = ~x_1379 & ~x_1380;
assign n_29141 = ~x_1381 & ~x_1382;
assign n_29142 =  n_29140 &  n_29141;
assign n_29143 =  n_29139 &  n_29142;
assign n_29144 =  n_29136 &  n_29143;
assign n_29145 = ~x_1359 & ~x_1360;
assign n_29146 = ~x_1361 & ~x_1362;
assign n_29147 =  n_29145 &  n_29146;
assign n_29148 = ~x_1355 & ~x_1356;
assign n_29149 = ~x_1357 & ~x_1358;
assign n_29150 =  n_29148 &  n_29149;
assign n_29151 =  n_29147 &  n_29150;
assign n_29152 = ~x_1367 & ~x_1368;
assign n_29153 = ~x_1369 & ~x_1370;
assign n_29154 =  n_29152 &  n_29153;
assign n_29155 = ~x_1363 & ~x_1364;
assign n_29156 = ~x_1365 & ~x_1366;
assign n_29157 =  n_29155 &  n_29156;
assign n_29158 =  n_29154 &  n_29157;
assign n_29159 =  n_29151 &  n_29158;
assign n_29160 =  n_29144 &  n_29159;
assign n_29161 =  n_28245 &  n_29160;
assign n_29162 = ~n_5192 & ~n_6531;
assign n_29163 = ~n_29161 &  n_29162;
assign n_29164 = ~n_28507 &  n_29163;
assign n_29165 = ~n_21107 & ~n_28508;
assign n_29166 =  n_3858 &  n_13015;
assign n_29167 = ~n_28859 & ~n_29166;
assign n_29168 =  n_29165 &  n_29167;
assign n_29169 =  n_29164 &  n_29168;
assign n_29170 =  n_3858 &  n_18433;
assign n_29171 =  n_27413 &  n_8254;
assign n_29172 = ~n_29171 & ~n_14817;
assign n_29173 = ~n_28728 & ~n_27911;
assign n_29174 =  n_29172 &  n_29173;
assign n_29175 = ~n_29170 &  n_29174;
assign n_29176 = ~n_13013 & ~n_24608;
assign n_29177 =  n_29176 &  n_28342;
assign n_29178 =  n_29175 &  n_29177;
assign n_29179 =  n_29169 &  n_29178;
assign n_29180 = ~n_28684 &  n_28828;
assign n_29181 =  n_585 &  n_27585;
assign n_29182 = ~n_29180 & ~n_29181;
assign n_29183 =  x_41 &  n_1180;
assign n_29184 = ~x_42 &  n_29183;
assign n_29185 = ~n_27637 &  n_27708;
assign n_29186 = ~n_29184 & ~n_29185;
assign n_29187 =  n_29182 &  n_29186;
assign n_29188 =  n_27424 &  n_1707;
assign n_29189 = ~n_8256 & ~n_10519;
assign n_29190 = ~n_29188 &  n_29189;
assign n_29191 =  n_29190 & ~n_13869;
assign n_29192 = ~n_27780 &  n_28350;
assign n_29193 =  n_28167 & ~n_28198;
assign n_29194 = ~n_29192 & ~n_29193;
assign n_29195 =  n_29191 &  n_29194;
assign n_29196 =  n_29187 &  n_29195;
assign n_29197 =  n_28535 &  n_3469;
assign n_29198 =  n_3858 &  n_28446;
assign n_29199 = ~n_29197 & ~n_29198;
assign n_29200 =  n_28240 &  n_3858;
assign n_29201 = ~n_22924 & ~n_29200;
assign n_29202 =  n_29199 &  n_29201;
assign n_29203 =  n_29202 & ~n_28019;
assign n_29204 =  n_29196 &  n_29203;
assign n_29205 =  n_29179 &  n_29204;
assign n_29206 =  n_29129 &  n_29205;
assign n_29207 =  n_29069 &  n_29206;
assign n_29208 =  n_29008 &  n_29207;
assign n_29209 =  n_29003 &  n_29208;
assign n_29210 = ~n_27426 &  n_29209;
assign n_29211 =  n_27254 &  n_28525;
assign n_29212 = ~n_29211 & ~n_27408;
assign n_29213 =  n_29210 &  n_29212;
assign n_29214 = ~n_28596 & ~n_27270;
assign n_29215 =  n_29213 &  n_29214;
assign n_29216 =  n_27399 &  n_28240;
assign n_29217 =  n_29216 &  n_2;
assign n_29218 = ~n_29217 & ~n_28570;
assign n_29219 =  n_27266 &  n_6530;
assign n_29220 =  n_27399 &  n_29219;
assign n_29221 = ~n_29220 & ~n_28579;
assign n_29222 =  n_27599 &  n_4993;
assign n_29223 =  n_29222 &  n_27399;
assign n_29224 =  n_27399 & ~n_28603;
assign n_29225 = ~n_29223 & ~n_29224;
assign n_29226 =  n_29221 &  n_29225;
assign n_29227 =  n_29218 &  n_29226;
assign n_29228 =  n_29215 &  n_29227;
assign n_29229 =  x_40 &  n_28609;
assign n_29230 =  n_19945 &  n_27273;
assign n_29231 =  n_27399 &  n_29230;
assign n_29232 = ~n_28564 & ~n_29231;
assign n_29233 = ~n_28617 &  n_29232;
assign n_29234 = ~n_29229 &  n_29233;
assign n_29235 =  n_28638 &  n_29234;
assign n_29236 =  n_29228 &  n_29235;
assign n_29237 =  n_28631 &  n_29236;
assign n_29238 =  n_26228 &  n_29237;
assign n_29239 =  x_40 & ~n_29238;
assign n_29240 = ~x_40 &  n_29238;
assign n_29241 = ~n_29239 & ~n_29240;
assign n_29242 = ~n_27599 & ~n_27268;
assign n_29243 =  n_3664 & ~n_29242;
assign n_29244 =  n_27399 &  n_28589;
assign n_29245 = ~n_27264 & ~n_29244;
assign n_29246 =  n_12420 &  n_27403;
assign n_29247 =  n_27399 &  n_29246;
assign n_29248 = ~n_28615 & ~n_29247;
assign n_29249 =  n_29245 &  n_29248;
assign n_29250 = ~n_29243 &  n_29249;
assign n_29251 = ~n_3276 & ~n_28715;
assign n_29252 =  n_1314 &  n_14808;
assign n_29253 =  n_29251 & ~n_29252;
assign n_29254 =  n_29253 & ~n_28694;
assign n_29255 =  n_4 &  n_28233;
assign n_29256 =  n_12420 &  n_29255;
assign n_29257 =  n_28131 &  n_29256;
assign n_29258 = ~n_28520 & ~n_29257;
assign n_29259 =  n_29254 &  n_29258;
assign n_29260 =  n_28319 &  n_28321;
assign n_29261 =  n_27258 &  n_784;
assign n_29262 = ~n_29261 & ~n_27598;
assign n_29263 = ~n_10517 &  n_29262;
assign n_29264 = ~n_29260 &  n_29263;
assign n_29265 = ~x_803 & ~x_804;
assign n_29266 = ~x_805 & ~x_806;
assign n_29267 =  n_29265 &  n_29266;
assign n_29268 = ~x_799 & ~x_800;
assign n_29269 = ~x_801 & ~x_802;
assign n_29270 =  n_29268 &  n_29269;
assign n_29271 =  n_29267 &  n_29270;
assign n_29272 = ~x_807 & ~x_808;
assign n_29273 = ~x_809 & ~x_810;
assign n_29274 =  n_29272 &  n_29273;
assign n_29275 =  n_4056 &  n_29274;
assign n_29276 =  n_29271 &  n_29275;
assign n_29277 = ~x_779 & ~x_780;
assign n_29278 = ~x_781 & ~x_782;
assign n_29279 =  n_29277 &  n_29278;
assign n_29280 =  n_5 &  n_29279;
assign n_29281 = ~x_787 & ~x_788;
assign n_29282 = ~x_789 & ~x_790;
assign n_29283 =  n_29281 &  n_29282;
assign n_29284 = ~x_783 & ~x_784;
assign n_29285 = ~x_785 & ~x_786;
assign n_29286 =  n_29284 &  n_29285;
assign n_29287 =  n_29283 &  n_29286;
assign n_29288 = ~x_795 & ~x_796;
assign n_29289 = ~x_797 & ~x_798;
assign n_29290 =  n_29288 &  n_29289;
assign n_29291 = ~x_791 & ~x_792;
assign n_29292 = ~x_793 & ~x_794;
assign n_29293 =  n_29291 &  n_29292;
assign n_29294 =  n_29290 &  n_29293;
assign n_29295 =  n_29287 &  n_29294;
assign n_29296 =  n_29280 &  n_29295;
assign n_29297 =  n_29276 &  n_29296;
assign n_29298 =  n_783 &  n_29297;
assign n_29299 = ~n_29298 & ~n_28019;
assign n_29300 =  n_29264 &  n_29299;
assign n_29301 =  n_29259 &  n_29300;
assign n_29302 =  n_29090 &  n_28870;
assign n_29303 =  n_28318 &  n_29302;
assign n_29304 = ~n_28533 & ~n_29084;
assign n_29305 =  n_29304 &  n_28854;
assign n_29306 =  n_29303 &  n_29305;
assign n_29307 =  n_28535 &  n_8254;
assign n_29308 =  n_29172 & ~n_29307;
assign n_29309 =  n_29308 &  n_28220;
assign n_29310 = ~n_27585 & ~n_13015;
assign n_29311 =  n_13014 & ~n_29310;
assign n_29312 = ~n_27782 & ~n_29311;
assign n_29313 =  n_29309 &  n_29312;
assign n_29314 =  n_29306 &  n_29313;
assign n_29315 =  n_28875 &  n_28431;
assign n_29316 =  n_28458 & ~n_27582;
assign n_29317 =  n_28864 & ~n_29316;
assign n_29318 =  n_29315 &  n_29317;
assign n_29319 = ~n_28230 &  n_29318;
assign n_29320 =  n_29314 &  n_29319;
assign n_29321 =  n_29301 &  n_29320;
assign n_29322 = ~n_27584 & ~n_27822;
assign n_29323 =  n_28929 &  n_29322;
assign n_29324 =  n_27669 &  n_27825;
assign n_29325 =  n_10518 &  n_27703;
assign n_29326 =  n_10318 &  n_29325;
assign n_29327 = ~n_29324 & ~n_29326;
assign n_29328 =  n_783 &  n_27406;
assign n_29329 = ~n_29328 & ~n_29122;
assign n_29330 = ~n_29170 & ~n_7866;
assign n_29331 = ~n_28467 & ~n_28199;
assign n_29332 =  n_29330 &  n_29331;
assign n_29333 =  n_29329 &  n_29332;
assign n_29334 =  n_29327 &  n_29333;
assign n_29335 =  n_27915 &  n_29334;
assign n_29336 =  n_29323 &  n_29335;
assign n_29337 =  n_29321 &  n_29336;
assign n_29338 =  n_28037 &  n_28441;
assign n_29339 = ~n_13667 & ~n_29338;
assign n_29340 =  n_29339 & ~n_8256;
assign n_29341 =  n_6533 &  n_3275;
assign n_29342 =  n_29340 & ~n_29341;
assign n_29343 =  n_783 &  n_6527;
assign n_29344 = ~n_29343 & ~n_4446;
assign n_29345 = ~n_12033 &  n_29344;
assign n_29346 =  n_28424 &  n_29345;
assign n_29347 = ~n_28846 &  n_29346;
assign n_29348 =  n_29342 &  n_29347;
assign n_29349 =  n_29006 &  n_28044;
assign n_29350 =  n_29348 &  n_29349;
assign n_29351 = ~n_29197 & ~n_28599;
assign n_29352 =  n_28331 &  n_29351;
assign n_29353 =  n_28535 &  n_783;
assign n_29354 = ~n_28914 & ~n_29353;
assign n_29355 = ~n_28866 &  n_29354;
assign n_29356 =  n_29352 &  n_29355;
assign n_29357 = ~n_1710 & ~n_13473;
assign n_29358 = ~n_28767 &  n_29357;
assign n_29359 = ~n_28324 &  n_29058;
assign n_29360 =  n_29358 &  n_29359;
assign n_29361 =  n_29356 &  n_29360;
assign n_29362 = ~n_27423 & ~n_27274;
assign n_29363 =  n_28115 & ~n_29362;
assign n_29364 = ~n_29363 & ~n_28823;
assign n_29365 = ~n_22345 &  n_28825;
assign n_29366 =  n_29364 &  n_29365;
assign n_29367 = ~n_20525 & ~n_29097;
assign n_29368 = ~n_6528 & ~n_28353;
assign n_29369 =  n_29367 &  n_29368;
assign n_29370 =  n_28391 & ~n_28422;
assign n_29371 = ~x_42 &  n_2304;
assign n_29372 = ~n_29370 & ~n_29371;
assign n_29373 =  n_29369 &  n_29372;
assign n_29374 =  n_29366 &  n_29373;
assign n_29375 =  n_29361 &  n_29374;
assign n_29376 = ~n_3665 & ~n_20332;
assign n_29377 = ~n_28829 & ~n_28511;
assign n_29378 =  n_29376 &  n_29377;
assign n_29379 = ~n_23503 & ~n_28727;
assign n_29380 =  n_28535 &  n_6533;
assign n_29381 = ~n_29380 & ~n_786;
assign n_29382 =  n_29379 &  n_29381;
assign n_29383 =  n_29378 &  n_29382;
assign n_29384 =  x_39 &  n_1;
assign n_29385 =  n_2499 &  n_29384;
assign n_29386 = ~n_28550 & ~n_29385;
assign n_29387 = ~n_28122 &  n_29386;
assign n_29388 = ~n_28778 & ~n_27588;
assign n_29389 = ~n_10519 & ~n_28723;
assign n_29390 = ~n_18448 &  n_29389;
assign n_29391 =  n_29388 &  n_29390;
assign n_29392 =  n_29387 &  n_29391;
assign n_29393 =  n_29383 &  n_29392;
assign n_29394 = ~n_28453 & ~n_28716;
assign n_29395 = ~n_28278 &  n_29394;
assign n_29396 =  n_783 &  n_27403;
assign n_29397 =  n_28336 & ~n_29396;
assign n_29398 =  n_29395 &  n_29397;
assign n_29399 = ~n_28644 & ~n_8824;
assign n_29400 = ~n_12421 &  n_29399;
assign n_29401 =  n_27266 &  n_783;
assign n_29402 = ~n_29401 & ~n_29064;
assign n_29403 = ~n_28722 & ~n_28436;
assign n_29404 =  n_29402 &  n_29403;
assign n_29405 =  n_29400 &  n_29404;
assign n_29406 = ~n_27596 & ~n_28523;
assign n_29407 =  n_29405 &  n_29406;
assign n_29408 =  n_29398 &  n_29407;
assign n_29409 =  n_29393 &  n_29408;
assign n_29410 =  n_29375 &  n_29409;
assign n_29411 =  n_28446 &  n_13014;
assign n_29412 = ~n_29411 & ~n_28461;
assign n_29413 = ~n_28214 & ~n_28987;
assign n_29414 =  n_29412 &  n_29413;
assign n_29415 =  n_27669 &  n_27670;
assign n_29416 =  n_29414 & ~n_29415;
assign n_29417 =  n_29011 &  n_29016;
assign n_29418 =  n_29416 &  n_29417;
assign n_29419 =  n_783 &  n_588;
assign n_29420 = ~n_29419 & ~n_28950;
assign n_29421 =  n_28530 &  n_29420;
assign n_29422 = ~n_27594 & ~n_28347;
assign n_29423 = ~n_6534 & ~n_5197;
assign n_29424 =  n_29422 &  n_29423;
assign n_29425 =  n_29421 &  n_29424;
assign n_29426 = ~n_28986 & ~n_28989;
assign n_29427 =  n_28446 &  n_12614;
assign n_29428 = ~n_29427 & ~n_28774;
assign n_29429 =  n_29426 &  n_29428;
assign n_29430 =  n_27923 &  n_28874;
assign n_29431 =  n_29429 &  n_29430;
assign n_29432 =  n_29425 &  n_29431;
assign n_29433 =  n_29418 &  n_29432;
assign n_29434 =  n_29410 &  n_29433;
assign n_29435 =  n_29350 &  n_29434;
assign n_29436 =  n_29337 &  n_29435;
assign n_29437 = ~n_28632 &  n_29436;
assign n_29438 = ~n_28617 &  n_29437;
assign n_29439 =  n_27262 &  n_979;
assign n_29440 = ~n_27254 &  n_29439;
assign n_29441 =  x_40 &  n_29440;
assign n_29442 =  n_27419 & ~n_29441;
assign n_29443 =  n_29438 &  n_29442;
assign n_29444 = ~n_27399 &  n_28602;
assign n_29445 = ~x_40 &  n_29440;
assign n_29446 = ~n_29444 & ~n_29445;
assign n_29447 =  n_27399 &  n_28578;
assign n_29448 =  x_40 &  n_28608;
assign n_29449 =  n_27399 &  n_29448;
assign n_29450 = ~n_27254 &  n_28586;
assign n_29451 = ~n_29449 & ~n_29450;
assign n_29452 = ~n_29447 &  n_29451;
assign n_29453 =  n_29446 &  n_29452;
assign n_29454 =  n_29443 &  n_29453;
assign n_29455 =  n_27399 &  n_27407;
assign n_29456 = ~n_28606 & ~n_29455;
assign n_29457 = ~n_28584 &  n_29456;
assign n_29458 = ~n_27254 &  n_27599;
assign n_29459 =  n_8818 &  n_29458;
assign n_29460 = ~n_29459 & ~n_28635;
assign n_29461 =  n_29457 &  n_29460;
assign n_29462 =  n_27399 &  n_28602;
assign n_29463 = ~n_27405 & ~n_28525;
assign n_29464 = ~n_29462 &  n_29463;
assign n_29465 =  n_29216 &  n_13012;
assign n_29466 = ~n_27261 & ~n_29465;
assign n_29467 =  n_29464 &  n_29466;
assign n_29468 =  n_29461 &  n_29467;
assign n_29469 =  n_29454 &  n_29468;
assign n_29470 =  n_29250 &  n_29469;
assign n_29471 = ~n_27129 &  n_29470;
assign n_29472 = ~n_28630 &  n_29471;
assign n_29473 =  n_25776 & ~n_26225;
assign n_29474 =  n_25320 & ~n_25772;
assign n_29475 = ~n_29473 & ~n_29474;
assign n_29476 =  n_29472 &  n_29475;
assign n_29477 =  x_39 & ~n_29476;
assign n_29478 = ~x_39 &  n_29476;
assign n_29479 = ~n_29477 & ~n_29478;
assign n_29480 =  n_29232 & ~n_27401;
assign n_29481 =  n_3664 &  n_29458;
assign n_29482 = ~n_29481 & ~n_27418;
assign n_29483 = ~n_28618 &  n_29482;
assign n_29484 =  n_29480 &  n_29483;
assign n_29485 =  n_28598 & ~n_29222;
assign n_29486 =  n_27599 &  n_12420;
assign n_29487 = ~n_29486 & ~n_27415;
assign n_29488 =  n_29485 &  n_29487;
assign n_29489 =  n_24413 & ~n_28037;
assign n_29490 = ~n_18445 & ~n_29489;
assign n_29491 =  n_1178 & ~n_29490;
assign n_29492 = ~n_29491 &  n_27714;
assign n_29493 =  n_27672 &  n_29492;
assign n_29494 =  n_29001 &  n_29493;
assign n_29495 =  n_28687 &  n_29323;
assign n_29496 =  n_29494 &  n_29495;
assign n_29497 = ~n_3663 & ~n_13002;
assign n_29498 =  n_1179 & ~n_29497;
assign n_29499 = ~n_8824 & ~n_29498;
assign n_29500 = ~n_28578 &  n_29499;
assign n_29501 = ~n_28547 &  n_29500;
assign n_29502 = ~n_29198 &  n_29114;
assign n_29503 =  n_29501 &  n_29502;
assign n_29504 = ~n_7479 & ~n_28770;
assign n_29505 =  n_28115 &  n_28758;
assign n_29506 = ~n_29505 & ~n_29419;
assign n_29507 =  n_29504 &  n_29506;
assign n_29508 = ~n_25775 & ~n_18446;
assign n_29509 = ~n_21686 & ~n_28126;
assign n_29510 =  n_29508 &  n_29509;
assign n_29511 = ~n_1907 & ~n_23698;
assign n_29512 =  n_29510 &  n_29511;
assign n_29513 =  n_29507 &  n_29512;
assign n_29514 =  n_29503 &  n_29513;
assign n_29515 = ~n_28467 & ~n_28781;
assign n_29516 = ~n_18448 & ~n_24414;
assign n_29517 =  n_29516 &  n_28203;
assign n_29518 =  n_29515 &  n_29517;
assign n_29519 = ~n_28863 & ~n_28279;
assign n_29520 = ~n_28447 &  n_29519;
assign n_29521 = ~x_895 & ~x_896;
assign n_29522 = ~x_897 & ~x_898;
assign n_29523 =  n_29521 &  n_29522;
assign n_29524 = ~x_891 & ~x_892;
assign n_29525 = ~x_893 & ~x_894;
assign n_29526 =  n_29524 &  n_29525;
assign n_29527 =  n_29523 &  n_29526;
assign n_29528 = ~x_903 & ~x_904;
assign n_29529 = ~x_905 & ~x_906;
assign n_29530 =  n_29528 &  n_29529;
assign n_29531 = ~x_899 & ~x_900;
assign n_29532 = ~x_901 & ~x_902;
assign n_29533 =  n_29531 &  n_29532;
assign n_29534 =  n_29530 &  n_29533;
assign n_29535 =  n_29527 &  n_29534;
assign n_29536 = ~x_879 & ~x_880;
assign n_29537 = ~x_881 & ~x_882;
assign n_29538 =  n_29536 &  n_29537;
assign n_29539 = ~x_875 & ~x_876;
assign n_29540 = ~x_877 & ~x_878;
assign n_29541 =  n_29539 &  n_29540;
assign n_29542 =  n_29538 &  n_29541;
assign n_29543 = ~x_887 & ~x_888;
assign n_29544 = ~x_889 & ~x_890;
assign n_29545 =  n_29543 &  n_29544;
assign n_29546 = ~x_883 & ~x_884;
assign n_29547 = ~x_885 & ~x_886;
assign n_29548 =  n_29546 &  n_29547;
assign n_29549 =  n_29545 &  n_29548;
assign n_29550 =  n_29542 &  n_29549;
assign n_29551 =  n_29535 &  n_29550;
assign n_29552 =  n_13014 &  n_13006;
assign n_29553 = ~n_29551 &  n_29552;
assign n_29554 = ~n_27586 & ~n_29553;
assign n_29555 =  n_29520 &  n_29554;
assign n_29556 =  n_29518 &  n_29555;
assign n_29557 =  n_29514 &  n_29556;
assign n_29558 = ~n_27596 & ~n_29080;
assign n_29559 =  n_29558 & ~n_29298;
assign n_29560 =  n_28245 & ~n_29160;
assign n_29561 = ~n_29560 & ~n_28278;
assign n_29562 =  n_29561 &  n_28339;
assign n_29563 =  n_29559 &  n_29562;
assign n_29564 = ~n_27924 & ~n_25776;
assign n_29565 = ~n_27840 & ~n_28165;
assign n_29566 =  n_29564 &  n_29565;
assign n_29567 = ~n_28716 & ~n_27601;
assign n_29568 = ~n_28114 & ~n_1710;
assign n_29569 =  n_29567 &  n_29568;
assign n_29570 =  n_29566 &  n_29569;
assign n_29571 =  n_2 &  n_6332;
assign n_29572 = ~n_29183 & ~n_29571;
assign n_29573 =  n_28745 &  n_29572;
assign n_29574 = ~n_28550 & ~n_10516;
assign n_29575 =  x_38 &  n_29401;
assign n_29576 = ~n_16334 & ~n_29575;
assign n_29577 =  n_29574 &  n_29576;
assign n_29578 =  n_29573 &  n_29577;
assign n_29579 =  n_29570 &  n_29578;
assign n_29580 =  n_29563 &  n_29579;
assign n_29581 =  n_29557 &  n_29580;
assign n_29582 =  n_29430 &  n_29414;
assign n_29583 =  n_29060 &  n_29582;
assign n_29584 =  n_28915 &  n_29054;
assign n_29585 = ~n_29584 &  n_29367;
assign n_29586 =  n_29368 &  n_28789;
assign n_29587 =  n_29585 &  n_29586;
assign n_29588 = ~n_27978 &  n_29587;
assign n_29589 = ~n_8808 & ~n_28706;
assign n_29590 = ~n_28426 &  n_29589;
assign n_29591 = ~n_28943 & ~n_29092;
assign n_29592 =  n_29590 &  n_29591;
assign n_29593 =  n_29592 &  n_28645;
assign n_29594 =  n_29588 &  n_29593;
assign n_29595 =  n_29583 &  n_29594;
assign n_29596 =  n_29581 &  n_29595;
assign n_29597 = ~n_3469 & ~n_13002;
assign n_29598 =  n_2499 & ~n_29597;
assign n_29599 =  n_28242 & ~n_29598;
assign n_29600 =  n_28318 &  n_29599;
assign n_29601 =  n_29600 &  n_27818;
assign n_29602 =  n_28458 &  n_27582;
assign n_29603 = ~n_29078 & ~n_28335;
assign n_29604 = ~n_3665 &  n_29603;
assign n_29605 = ~n_29602 &  n_29604;
assign n_29606 =  n_29605 &  n_29340;
assign n_29607 =  n_29601 &  n_29606;
assign n_29608 = ~x_40 &  n_28754;
assign n_29609 = ~n_12809 & ~n_29608;
assign n_29610 = ~n_3276 & ~n_12421;
assign n_29611 = ~n_21879 &  n_29610;
assign n_29612 = ~n_12616 &  n_29611;
assign n_29613 =  n_29609 &  n_29612;
assign n_29614 =  n_28983 &  n_29613;
assign n_29615 = ~n_28390 & ~n_28722;
assign n_29616 =  n_27406 & ~n_23897;
assign n_29617 = ~n_29616 & ~n_29161;
assign n_29618 =  n_29615 &  n_29617;
assign n_29619 =  n_27595 &  n_29329;
assign n_29620 =  n_29618 &  n_29619;
assign n_29621 =  n_29614 &  n_29620;
assign n_29622 =  n_24801 &  n_27403;
assign n_29623 =  n_3664 &  n_6527;
assign n_29624 = ~n_29623 & ~n_28326;
assign n_29625 = ~n_29622 &  n_29624;
assign n_29626 = ~x_42 &  n_13868;
assign n_29627 = ~n_29070 & ~n_29626;
assign n_29628 =  n_29625 &  n_29627;
assign n_29629 =  n_28735 &  n_29628;
assign n_29630 = ~n_14812 &  n_28740;
assign n_29631 =  n_29175 &  n_29630;
assign n_29632 =  n_29629 &  n_29631;
assign n_29633 =  n_29621 &  n_29632;
assign n_29634 =  n_29607 &  n_29633;
assign n_29635 =  n_29596 &  n_29634;
assign n_29636 =  n_10319 &  n_188;
assign n_29637 =  n_12614 &  n_29636;
assign n_29638 =  n_28232 &  n_29637;
assign n_29639 = ~n_29638 & ~n_28133;
assign n_29640 =  n_1708 &  n_28022;
assign n_29641 = ~n_29343 & ~n_29640;
assign n_29642 =  n_29258 &  n_29641;
assign n_29643 =  n_29639 &  n_29642;
assign n_29644 =  n_28237 &  n_29643;
assign n_29645 =  n_13014 &  n_29325;
assign n_29646 =  n_27582 &  n_27583;
assign n_29647 = ~n_27836 & ~n_29646;
assign n_29648 = ~n_29645 &  n_29647;
assign n_29649 = ~n_28119 &  n_29648;
assign n_29650 = ~n_28024 &  n_29649;
assign n_29651 =  n_28642 &  n_29650;
assign n_29652 =  n_29644 &  n_29651;
assign n_29653 =  n_29635 &  n_29652;
assign n_29654 =  n_29496 &  n_29653;
assign n_29655 = ~n_28571 &  n_29654;
assign n_29656 = ~n_28587 &  n_29655;
assign n_29657 =  n_8060 &  n_27403;
assign n_29658 =  n_27399 &  n_29657;
assign n_29659 = ~n_28567 & ~n_29658;
assign n_29660 =  n_29659 & ~n_28615;
assign n_29661 =  n_29656 &  n_29660;
assign n_29662 =  n_29488 &  n_29661;
assign n_29663 =  n_29484 &  n_29662;
assign n_29664 = ~n_27129 &  n_29663;
assign n_29665 =  x_38 & ~n_29664;
assign n_29666 = ~x_38 &  n_29664;
assign n_29667 = ~n_29665 & ~n_29666;
assign n_29668 = ~x_1000 & ~x_1001;
assign n_29669 = ~x_999 &  n_29668;
assign n_29670 = ~x_998 &  n_29669;
assign n_29671 = ~x_997 & ~x_1002;
assign n_29672 =  n_29670 &  n_29671;
assign n_29673 = ~x_996 &  n_29672;
assign n_29674 = ~x_995 &  n_29673;
assign n_29675 = ~x_994 &  n_29674;
assign n_29676 = ~x_993 &  n_29675;
assign n_29677 = ~x_992 &  n_29676;
assign n_29678 = ~x_991 &  n_29677;
assign n_29679 = ~x_990 &  n_29678;
assign n_29680 = ~x_989 &  n_29679;
assign n_29681 = ~x_988 &  n_29680;
assign n_29682 = ~x_987 &  n_29681;
assign n_29683 = ~x_986 &  n_29682;
assign n_29684 = ~x_985 &  n_29683;
assign n_29685 = ~x_984 &  n_29684;
assign n_29686 = ~x_983 &  n_29685;
assign n_29687 = ~x_982 &  n_29686;
assign n_29688 = ~x_981 &  n_29687;
assign n_29689 = ~x_980 &  n_29688;
assign n_29690 = ~x_979 &  n_29689;
assign n_29691 = ~x_978 &  n_29690;
assign n_29692 = ~x_977 &  n_29691;
assign n_29693 = ~x_976 &  n_29692;
assign n_29694 = ~x_975 &  n_29693;
assign n_29695 = ~x_974 &  n_29694;
assign n_29696 = ~x_973 &  n_29695;
assign n_29697 =  x_973 & ~n_29695;
assign n_29698 = ~n_29696 & ~n_29697;
assign n_29699 =  x_975 & ~n_29693;
assign n_29700 = ~n_29694 & ~n_29699;
assign n_29701 =  x_977 & ~n_29691;
assign n_29702 = ~n_29692 & ~n_29701;
assign n_29703 =  x_979 & ~n_29689;
assign n_29704 = ~n_29690 & ~n_29703;
assign n_29705 =  x_981 & ~n_29687;
assign n_29706 = ~n_29688 & ~n_29705;
assign n_29707 =  x_983 & ~n_29685;
assign n_29708 = ~n_29686 & ~n_29707;
assign n_29709 =  x_985 & ~n_29683;
assign n_29710 = ~n_29684 & ~n_29709;
assign n_29711 =  x_987 & ~n_29681;
assign n_29712 = ~n_29682 & ~n_29711;
assign n_29713 =  x_989 & ~n_29679;
assign n_29714 = ~n_29680 & ~n_29713;
assign n_29715 =  x_991 & ~n_29677;
assign n_29716 = ~n_29678 & ~n_29715;
assign n_29717 =  x_993 & ~n_29675;
assign n_29718 = ~n_29676 & ~n_29717;
assign n_29719 =  x_995 & ~n_29673;
assign n_29720 = ~n_29674 & ~n_29719;
assign n_29721 = ~x_997 &  x_1002;
assign n_29722 =  n_29670 &  n_29721;
assign n_29723 = ~x_996 &  n_29722;
assign n_29724 =  n_29720 &  n_29723;
assign n_29725 = ~x_994 &  n_29724;
assign n_29726 =  n_29718 &  n_29725;
assign n_29727 = ~x_992 &  n_29726;
assign n_29728 =  n_29716 &  n_29727;
assign n_29729 = ~x_990 &  n_29728;
assign n_29730 =  n_29714 &  n_29729;
assign n_29731 = ~x_988 &  n_29730;
assign n_29732 =  n_29712 &  n_29731;
assign n_29733 = ~x_986 &  n_29732;
assign n_29734 =  n_29710 &  n_29733;
assign n_29735 = ~x_984 &  n_29734;
assign n_29736 =  n_29708 &  n_29735;
assign n_29737 = ~x_982 &  n_29736;
assign n_29738 =  n_29706 &  n_29737;
assign n_29739 = ~x_980 &  n_29738;
assign n_29740 =  n_29704 &  n_29739;
assign n_29741 = ~x_978 &  n_29740;
assign n_29742 =  n_29702 &  n_29741;
assign n_29743 = ~x_976 &  n_29742;
assign n_29744 =  n_29700 &  n_29743;
assign n_29745 = ~x_974 &  n_29744;
assign n_29746 =  n_29698 &  n_29745;
assign n_29747 = ~x_972 &  n_29746;
assign n_29748 = ~x_972 &  n_29696;
assign n_29749 = ~x_971 & ~n_29748;
assign n_29750 =  x_971 &  n_29748;
assign n_29751 = ~n_29749 & ~n_29750;
assign n_29752 = ~n_29747 &  n_29751;
assign n_29753 =  n_29747 & ~n_29751;
assign n_29754 = ~n_29752 & ~n_29753;
assign n_29755 =  x_972 & ~n_29696;
assign n_29756 = ~n_29748 & ~n_29755;
assign n_29757 = ~n_29746 & ~n_29756;
assign n_29758 = ~n_29747 & ~n_29757;
assign n_29759 = ~n_29698 & ~n_29745;
assign n_29760 = ~n_29746 & ~n_29759;
assign n_29761 =  x_974 & ~n_29694;
assign n_29762 = ~n_29695 & ~n_29761;
assign n_29763 = ~n_29744 & ~n_29762;
assign n_29764 = ~n_29745 & ~n_29763;
assign n_29765 = ~n_29700 & ~n_29743;
assign n_29766 = ~n_29744 & ~n_29765;
assign n_29767 =  x_976 & ~n_29692;
assign n_29768 = ~n_29693 & ~n_29767;
assign n_29769 = ~n_29742 & ~n_29768;
assign n_29770 = ~n_29743 & ~n_29769;
assign n_29771 = ~n_29702 & ~n_29741;
assign n_29772 = ~n_29742 & ~n_29771;
assign n_29773 =  x_978 & ~n_29690;
assign n_29774 = ~n_29691 & ~n_29773;
assign n_29775 = ~n_29740 & ~n_29774;
assign n_29776 = ~n_29741 & ~n_29775;
assign n_29777 = ~n_29704 & ~n_29739;
assign n_29778 = ~n_29740 & ~n_29777;
assign n_29779 =  x_980 & ~n_29688;
assign n_29780 = ~n_29689 & ~n_29779;
assign n_29781 = ~n_29738 & ~n_29780;
assign n_29782 = ~n_29739 & ~n_29781;
assign n_29783 = ~n_29706 & ~n_29737;
assign n_29784 = ~n_29738 & ~n_29783;
assign n_29785 =  x_982 & ~n_29686;
assign n_29786 = ~n_29687 & ~n_29785;
assign n_29787 = ~n_29736 & ~n_29786;
assign n_29788 = ~n_29737 & ~n_29787;
assign n_29789 = ~n_29708 & ~n_29735;
assign n_29790 = ~n_29736 & ~n_29789;
assign n_29791 =  x_984 & ~n_29684;
assign n_29792 = ~n_29685 & ~n_29791;
assign n_29793 = ~n_29734 & ~n_29792;
assign n_29794 = ~n_29735 & ~n_29793;
assign n_29795 = ~n_29710 & ~n_29733;
assign n_29796 = ~n_29734 & ~n_29795;
assign n_29797 =  x_986 & ~n_29682;
assign n_29798 = ~n_29683 & ~n_29797;
assign n_29799 = ~n_29732 & ~n_29798;
assign n_29800 = ~n_29733 & ~n_29799;
assign n_29801 = ~n_29712 & ~n_29731;
assign n_29802 = ~n_29732 & ~n_29801;
assign n_29803 =  x_988 & ~n_29680;
assign n_29804 = ~n_29681 & ~n_29803;
assign n_29805 = ~n_29730 & ~n_29804;
assign n_29806 = ~n_29731 & ~n_29805;
assign n_29807 = ~n_29714 & ~n_29729;
assign n_29808 = ~n_29730 & ~n_29807;
assign n_29809 =  x_990 & ~n_29678;
assign n_29810 = ~n_29679 & ~n_29809;
assign n_29811 = ~n_29728 & ~n_29810;
assign n_29812 = ~n_29729 & ~n_29811;
assign n_29813 = ~n_29716 & ~n_29727;
assign n_29814 = ~n_29728 & ~n_29813;
assign n_29815 =  x_992 & ~n_29676;
assign n_29816 = ~n_29677 & ~n_29815;
assign n_29817 = ~n_29726 & ~n_29816;
assign n_29818 = ~n_29727 & ~n_29817;
assign n_29819 = ~n_29718 & ~n_29725;
assign n_29820 = ~n_29726 & ~n_29819;
assign n_29821 =  x_994 & ~n_29674;
assign n_29822 = ~n_29675 & ~n_29821;
assign n_29823 = ~n_29724 & ~n_29822;
assign n_29824 = ~n_29725 & ~n_29823;
assign n_29825 = ~n_29720 & ~n_29723;
assign n_29826 = ~n_29724 & ~n_29825;
assign n_29827 = ~n_29672 & ~n_29722;
assign n_29828 =  x_996 & ~n_29827;
assign n_29829 = ~x_996 &  n_29827;
assign n_29830 = ~n_29828 & ~n_29829;
assign n_29831 =  x_997 & ~n_29670;
assign n_29832 =  n_29827 & ~n_29831;
assign n_29833 =  x_999 & ~n_29668;
assign n_29834 = ~n_29669 & ~n_29833;
assign n_29835 = ~x_969 & ~x_1001;
assign n_29836 =  x_970 & ~x_1002;
assign n_29837 =  x_969 &  x_1001;
assign n_29838 = ~n_29836 & ~n_29837;
assign n_29839 = ~n_29835 & ~n_29838;
assign n_29840 = ~x_968 & ~n_29839;
assign n_29841 =  x_1000 & ~x_1001;
assign n_29842 = ~x_1000 &  x_1001;
assign n_29843 = ~n_29841 & ~n_29842;
assign n_29844 =  x_968 &  n_29839;
assign n_29845 =  n_29843 & ~n_29844;
assign n_29846 = ~n_29840 & ~n_29845;
assign n_29847 = ~n_29834 & ~n_29846;
assign n_29848 =  n_29834 &  n_29846;
assign n_29849 = ~x_967 & ~n_29848;
assign n_29850 = ~n_29847 & ~n_29849;
assign n_29851 =  x_998 & ~n_29669;
assign n_29852 = ~n_29670 & ~n_29851;
assign n_29853 = ~n_29850 & ~n_29852;
assign n_29854 =  n_29850 &  n_29852;
assign n_29855 = ~x_966 & ~n_29854;
assign n_29856 = ~n_29853 & ~n_29855;
assign n_29857 = ~n_29832 & ~n_29856;
assign n_29858 =  n_29832 &  n_29856;
assign n_29859 = ~x_965 & ~n_29858;
assign n_29860 = ~n_29857 & ~n_29859;
assign n_29861 =  n_29830 & ~n_29860;
assign n_29862 = ~n_29830 &  n_29860;
assign n_29863 = ~x_964 & ~n_29862;
assign n_29864 = ~n_29861 & ~n_29863;
assign n_29865 = ~n_29826 & ~n_29864;
assign n_29866 =  n_29826 &  n_29864;
assign n_29867 = ~x_963 & ~n_29866;
assign n_29868 = ~n_29865 & ~n_29867;
assign n_29869 = ~n_29824 & ~n_29868;
assign n_29870 =  n_29824 &  n_29868;
assign n_29871 = ~x_962 & ~n_29870;
assign n_29872 = ~n_29869 & ~n_29871;
assign n_29873 = ~n_29820 & ~n_29872;
assign n_29874 =  n_29820 &  n_29872;
assign n_29875 = ~x_961 & ~n_29874;
assign n_29876 = ~n_29873 & ~n_29875;
assign n_29877 = ~n_29818 & ~n_29876;
assign n_29878 =  n_29818 &  n_29876;
assign n_29879 = ~x_960 & ~n_29878;
assign n_29880 = ~n_29877 & ~n_29879;
assign n_29881 = ~n_29814 & ~n_29880;
assign n_29882 =  n_29814 &  n_29880;
assign n_29883 = ~x_959 & ~n_29882;
assign n_29884 = ~n_29881 & ~n_29883;
assign n_29885 = ~n_29812 & ~n_29884;
assign n_29886 =  n_29812 &  n_29884;
assign n_29887 = ~x_958 & ~n_29886;
assign n_29888 = ~n_29885 & ~n_29887;
assign n_29889 = ~n_29808 & ~n_29888;
assign n_29890 =  n_29808 &  n_29888;
assign n_29891 = ~x_957 & ~n_29890;
assign n_29892 = ~n_29889 & ~n_29891;
assign n_29893 = ~n_29806 & ~n_29892;
assign n_29894 =  n_29806 &  n_29892;
assign n_29895 = ~x_956 & ~n_29894;
assign n_29896 = ~n_29893 & ~n_29895;
assign n_29897 = ~n_29802 & ~n_29896;
assign n_29898 =  n_29802 &  n_29896;
assign n_29899 = ~x_955 & ~n_29898;
assign n_29900 = ~n_29897 & ~n_29899;
assign n_29901 = ~n_29800 & ~n_29900;
assign n_29902 =  n_29800 &  n_29900;
assign n_29903 = ~x_954 & ~n_29902;
assign n_29904 = ~n_29901 & ~n_29903;
assign n_29905 = ~n_29796 & ~n_29904;
assign n_29906 =  n_29796 &  n_29904;
assign n_29907 = ~x_953 & ~n_29906;
assign n_29908 = ~n_29905 & ~n_29907;
assign n_29909 = ~n_29794 & ~n_29908;
assign n_29910 =  n_29794 &  n_29908;
assign n_29911 = ~x_952 & ~n_29910;
assign n_29912 = ~n_29909 & ~n_29911;
assign n_29913 = ~n_29790 & ~n_29912;
assign n_29914 =  n_29790 &  n_29912;
assign n_29915 = ~x_951 & ~n_29914;
assign n_29916 = ~n_29913 & ~n_29915;
assign n_29917 = ~n_29788 & ~n_29916;
assign n_29918 =  n_29788 &  n_29916;
assign n_29919 = ~x_950 & ~n_29918;
assign n_29920 = ~n_29917 & ~n_29919;
assign n_29921 = ~n_29784 & ~n_29920;
assign n_29922 =  n_29784 &  n_29920;
assign n_29923 = ~x_949 & ~n_29922;
assign n_29924 = ~n_29921 & ~n_29923;
assign n_29925 = ~n_29782 & ~n_29924;
assign n_29926 =  n_29782 &  n_29924;
assign n_29927 = ~x_948 & ~n_29926;
assign n_29928 = ~n_29925 & ~n_29927;
assign n_29929 = ~n_29778 & ~n_29928;
assign n_29930 =  n_29778 &  n_29928;
assign n_29931 = ~x_947 & ~n_29930;
assign n_29932 = ~n_29929 & ~n_29931;
assign n_29933 = ~n_29776 & ~n_29932;
assign n_29934 =  n_29776 &  n_29932;
assign n_29935 = ~x_946 & ~n_29934;
assign n_29936 = ~n_29933 & ~n_29935;
assign n_29937 = ~n_29772 & ~n_29936;
assign n_29938 =  n_29772 &  n_29936;
assign n_29939 = ~x_945 & ~n_29938;
assign n_29940 = ~n_29937 & ~n_29939;
assign n_29941 = ~n_29770 & ~n_29940;
assign n_29942 =  n_29770 &  n_29940;
assign n_29943 = ~x_944 & ~n_29942;
assign n_29944 = ~n_29941 & ~n_29943;
assign n_29945 = ~n_29766 & ~n_29944;
assign n_29946 =  n_29766 &  n_29944;
assign n_29947 = ~x_943 & ~n_29946;
assign n_29948 = ~n_29945 & ~n_29947;
assign n_29949 = ~n_29764 & ~n_29948;
assign n_29950 =  n_29764 &  n_29948;
assign n_29951 = ~x_942 & ~n_29950;
assign n_29952 = ~n_29949 & ~n_29951;
assign n_29953 = ~n_29760 & ~n_29952;
assign n_29954 =  n_29760 &  n_29952;
assign n_29955 = ~x_941 & ~n_29954;
assign n_29956 = ~n_29953 & ~n_29955;
assign n_29957 = ~n_29758 & ~n_29956;
assign n_29958 =  n_29758 &  n_29956;
assign n_29959 = ~x_940 & ~n_29958;
assign n_29960 = ~n_29957 & ~n_29959;
assign n_29961 =  n_29754 &  n_29960;
assign n_29962 = ~n_29754 & ~n_29960;
assign n_29963 = ~n_29961 & ~n_29962;
assign n_29964 = ~x_939 & ~n_29963;
assign n_29965 =  x_939 &  n_29963;
assign n_29966 = ~n_29964 & ~n_29965;
assign n_29967 = ~n_29957 & ~n_29958;
assign n_29968 =  x_940 &  n_29967;
assign n_29969 = ~x_940 & ~n_29967;
assign n_29970 = ~n_29968 & ~n_29969;
assign n_29971 = ~n_29747 &  n_29749;
assign n_29972 = ~n_29960 &  n_29971;
assign n_29973 = ~n_29953 & ~n_29954;
assign n_29974 =  x_941 &  n_29973;
assign n_29975 = ~x_941 & ~n_29973;
assign n_29976 = ~n_29974 & ~n_29975;
assign n_29977 = ~n_29949 & ~n_29950;
assign n_29978 =  x_942 &  n_29977;
assign n_29979 = ~x_942 & ~n_29977;
assign n_29980 = ~n_29978 & ~n_29979;
assign n_29981 = ~n_29945 & ~n_29946;
assign n_29982 =  x_943 &  n_29981;
assign n_29983 = ~x_943 & ~n_29981;
assign n_29984 = ~n_29982 & ~n_29983;
assign n_29985 = ~n_29941 & ~n_29942;
assign n_29986 =  x_944 &  n_29985;
assign n_29987 = ~x_944 & ~n_29985;
assign n_29988 = ~n_29986 & ~n_29987;
assign n_29989 = ~n_29937 & ~n_29938;
assign n_29990 =  x_945 &  n_29989;
assign n_29991 = ~x_945 & ~n_29989;
assign n_29992 = ~n_29990 & ~n_29991;
assign n_29993 = ~n_29933 & ~n_29934;
assign n_29994 =  x_946 &  n_29993;
assign n_29995 = ~x_946 & ~n_29993;
assign n_29996 = ~n_29994 & ~n_29995;
assign n_29997 = ~n_29929 & ~n_29930;
assign n_29998 =  x_947 &  n_29997;
assign n_29999 = ~x_947 & ~n_29997;
assign n_30000 = ~n_29998 & ~n_29999;
assign n_30001 = ~n_29925 & ~n_29926;
assign n_30002 =  x_948 &  n_30001;
assign n_30003 = ~x_948 & ~n_30001;
assign n_30004 = ~n_30002 & ~n_30003;
assign n_30005 = ~n_29921 & ~n_29922;
assign n_30006 =  x_949 &  n_30005;
assign n_30007 = ~x_949 & ~n_30005;
assign n_30008 = ~n_30006 & ~n_30007;
assign n_30009 = ~n_29917 & ~n_29918;
assign n_30010 =  x_950 &  n_30009;
assign n_30011 = ~x_950 & ~n_30009;
assign n_30012 = ~n_30010 & ~n_30011;
assign n_30013 = ~n_29913 & ~n_29914;
assign n_30014 =  x_951 &  n_30013;
assign n_30015 = ~x_951 & ~n_30013;
assign n_30016 = ~n_30014 & ~n_30015;
assign n_30017 = ~n_29909 & ~n_29910;
assign n_30018 =  x_952 &  n_30017;
assign n_30019 = ~x_952 & ~n_30017;
assign n_30020 = ~n_30018 & ~n_30019;
assign n_30021 = ~n_29905 & ~n_29906;
assign n_30022 =  x_953 &  n_30021;
assign n_30023 = ~x_953 & ~n_30021;
assign n_30024 = ~n_30022 & ~n_30023;
assign n_30025 = ~n_29901 & ~n_29902;
assign n_30026 =  x_954 &  n_30025;
assign n_30027 = ~x_954 & ~n_30025;
assign n_30028 = ~n_30026 & ~n_30027;
assign n_30029 = ~n_29897 & ~n_29898;
assign n_30030 =  x_955 &  n_30029;
assign n_30031 = ~x_955 & ~n_30029;
assign n_30032 = ~n_30030 & ~n_30031;
assign n_30033 = ~n_29893 & ~n_29894;
assign n_30034 =  x_956 &  n_30033;
assign n_30035 = ~x_956 & ~n_30033;
assign n_30036 = ~n_30034 & ~n_30035;
assign n_30037 = ~n_29889 & ~n_29890;
assign n_30038 =  x_957 &  n_30037;
assign n_30039 = ~x_957 & ~n_30037;
assign n_30040 = ~n_30038 & ~n_30039;
assign n_30041 = ~n_29885 & ~n_29886;
assign n_30042 =  x_958 &  n_30041;
assign n_30043 = ~x_958 & ~n_30041;
assign n_30044 = ~n_30042 & ~n_30043;
assign n_30045 = ~n_29881 & ~n_29882;
assign n_30046 =  x_959 &  n_30045;
assign n_30047 = ~x_959 & ~n_30045;
assign n_30048 = ~n_30046 & ~n_30047;
assign n_30049 = ~n_29877 & ~n_29878;
assign n_30050 =  x_960 &  n_30049;
assign n_30051 = ~x_960 & ~n_30049;
assign n_30052 = ~n_30050 & ~n_30051;
assign n_30053 = ~n_29873 & ~n_29874;
assign n_30054 =  x_961 &  n_30053;
assign n_30055 = ~x_961 & ~n_30053;
assign n_30056 = ~n_30054 & ~n_30055;
assign n_30057 = ~n_29869 & ~n_29870;
assign n_30058 =  x_962 &  n_30057;
assign n_30059 = ~x_962 & ~n_30057;
assign n_30060 = ~n_30058 & ~n_30059;
assign n_30061 = ~n_29865 & ~n_29866;
assign n_30062 =  x_963 &  n_30061;
assign n_30063 = ~x_963 & ~n_30061;
assign n_30064 = ~n_30062 & ~n_30063;
assign n_30065 = ~n_29861 & ~n_29862;
assign n_30066 =  x_964 &  n_30065;
assign n_30067 = ~x_964 & ~n_30065;
assign n_30068 = ~n_30066 & ~n_30067;
assign n_30069 = ~n_29857 & ~n_29858;
assign n_30070 =  x_965 &  n_30069;
assign n_30071 = ~x_965 & ~n_30069;
assign n_30072 = ~n_30070 & ~n_30071;
assign n_30073 = ~n_29853 & ~n_29854;
assign n_30074 =  x_966 &  n_30073;
assign n_30075 = ~x_966 & ~n_30073;
assign n_30076 = ~n_30074 & ~n_30075;
assign n_30077 = ~n_29847 & ~n_29848;
assign n_30078 =  x_967 &  n_30077;
assign n_30079 = ~x_967 & ~n_30077;
assign n_30080 = ~n_30078 & ~n_30079;
assign n_30081 = ~n_29840 & ~n_29844;
assign n_30082 = ~n_29843 & ~n_30081;
assign n_30083 = ~n_29840 &  n_29845;
assign n_30084 = ~n_29835 & ~n_29837;
assign n_30085 = ~x_970 &  x_1002;
assign n_30086 = ~n_29836 & ~n_30085;
assign n_30087 = ~n_30084 &  n_30086;
assign n_30088 = ~n_30083 &  n_30087;
assign n_30089 = ~n_30082 &  n_30088;
assign n_30090 = ~n_30080 &  n_30089;
assign n_30091 = ~n_30076 &  n_30090;
assign n_30092 = ~n_30072 &  n_30091;
assign n_30093 = ~n_30068 &  n_30092;
assign n_30094 = ~n_30064 &  n_30093;
assign n_30095 = ~n_30060 &  n_30094;
assign n_30096 = ~n_30056 &  n_30095;
assign n_30097 = ~n_30052 &  n_30096;
assign n_30098 = ~n_30048 &  n_30097;
assign n_30099 = ~n_30044 &  n_30098;
assign n_30100 = ~n_30040 &  n_30099;
assign n_30101 = ~n_30036 &  n_30100;
assign n_30102 = ~n_30032 &  n_30101;
assign n_30103 = ~n_30028 &  n_30102;
assign n_30104 = ~n_30024 &  n_30103;
assign n_30105 = ~n_30020 &  n_30104;
assign n_30106 = ~n_30016 &  n_30105;
assign n_30107 = ~n_30012 &  n_30106;
assign n_30108 = ~n_30008 &  n_30107;
assign n_30109 = ~n_30004 &  n_30108;
assign n_30110 = ~n_30000 &  n_30109;
assign n_30111 = ~n_29996 &  n_30110;
assign n_30112 = ~n_29992 &  n_30111;
assign n_30113 = ~n_29988 &  n_30112;
assign n_30114 = ~n_29984 &  n_30113;
assign n_30115 = ~n_29980 &  n_30114;
assign n_30116 = ~n_29976 &  n_30115;
assign n_30117 = ~n_29972 &  n_30116;
assign n_30118 = ~n_29970 &  n_30117;
assign n_30119 = ~n_29966 &  n_30118;
assign n_30120 =  n_28550 &  n_30119;
assign n_30121 = ~x_1896 & ~x_1897;
assign n_30122 = ~x_1895 &  n_30121;
assign n_30123 = ~x_1894 &  n_30122;
assign n_30124 = ~x_1893 & ~x_1898;
assign n_30125 =  n_30123 &  n_30124;
assign n_30126 = ~x_1892 &  n_30125;
assign n_30127 = ~x_1891 &  n_30126;
assign n_30128 = ~x_1890 &  n_30127;
assign n_30129 = ~x_1889 &  n_30128;
assign n_30130 = ~x_1888 &  n_30129;
assign n_30131 = ~x_1887 &  n_30130;
assign n_30132 = ~x_1886 &  n_30131;
assign n_30133 = ~x_1885 &  n_30132;
assign n_30134 = ~x_1884 &  n_30133;
assign n_30135 = ~x_1883 &  n_30134;
assign n_30136 = ~x_1882 &  n_30135;
assign n_30137 = ~x_1881 &  n_30136;
assign n_30138 = ~x_1880 &  n_30137;
assign n_30139 = ~x_1879 &  n_30138;
assign n_30140 = ~x_1878 &  n_30139;
assign n_30141 = ~x_1877 &  n_30140;
assign n_30142 = ~x_1876 &  n_30141;
assign n_30143 = ~x_1875 &  n_30142;
assign n_30144 = ~x_1874 &  n_30143;
assign n_30145 = ~x_1873 &  n_30144;
assign n_30146 = ~x_1872 &  n_30145;
assign n_30147 = ~x_1871 &  n_30146;
assign n_30148 =  x_1871 & ~n_30146;
assign n_30149 = ~n_30147 & ~n_30148;
assign n_30150 =  x_1873 & ~n_30144;
assign n_30151 = ~n_30145 & ~n_30150;
assign n_30152 =  x_1875 & ~n_30142;
assign n_30153 = ~n_30143 & ~n_30152;
assign n_30154 =  x_1877 & ~n_30140;
assign n_30155 = ~n_30141 & ~n_30154;
assign n_30156 =  x_1879 & ~n_30138;
assign n_30157 = ~n_30139 & ~n_30156;
assign n_30158 =  x_1881 & ~n_30136;
assign n_30159 = ~n_30137 & ~n_30158;
assign n_30160 =  x_1883 & ~n_30134;
assign n_30161 = ~n_30135 & ~n_30160;
assign n_30162 =  x_1885 & ~n_30132;
assign n_30163 = ~n_30133 & ~n_30162;
assign n_30164 =  x_1887 & ~n_30130;
assign n_30165 = ~n_30131 & ~n_30164;
assign n_30166 =  x_1889 & ~n_30128;
assign n_30167 = ~n_30129 & ~n_30166;
assign n_30168 =  x_1891 & ~n_30126;
assign n_30169 = ~n_30127 & ~n_30168;
assign n_30170 = ~x_1893 &  x_1898;
assign n_30171 =  n_30123 &  n_30170;
assign n_30172 = ~x_1892 &  n_30171;
assign n_30173 =  n_30169 &  n_30172;
assign n_30174 = ~x_1890 &  n_30173;
assign n_30175 =  n_30167 &  n_30174;
assign n_30176 = ~x_1888 &  n_30175;
assign n_30177 =  n_30165 &  n_30176;
assign n_30178 = ~x_1886 &  n_30177;
assign n_30179 =  n_30163 &  n_30178;
assign n_30180 = ~x_1884 &  n_30179;
assign n_30181 =  n_30161 &  n_30180;
assign n_30182 = ~x_1882 &  n_30181;
assign n_30183 =  n_30159 &  n_30182;
assign n_30184 = ~x_1880 &  n_30183;
assign n_30185 =  n_30157 &  n_30184;
assign n_30186 = ~x_1878 &  n_30185;
assign n_30187 =  n_30155 &  n_30186;
assign n_30188 = ~x_1876 &  n_30187;
assign n_30189 =  n_30153 &  n_30188;
assign n_30190 = ~x_1874 &  n_30189;
assign n_30191 =  n_30151 &  n_30190;
assign n_30192 = ~x_1872 &  n_30191;
assign n_30193 =  n_30149 &  n_30192;
assign n_30194 = ~x_1870 &  n_30193;
assign n_30195 = ~x_1870 &  n_30147;
assign n_30196 = ~x_1869 &  n_30195;
assign n_30197 =  x_1869 & ~n_30195;
assign n_30198 = ~n_30196 & ~n_30197;
assign n_30199 =  n_30194 &  n_30198;
assign n_30200 = ~x_1868 &  n_30199;
assign n_30201 = ~x_1868 &  n_30196;
assign n_30202 =  x_1868 & ~n_30196;
assign n_30203 = ~n_30201 & ~n_30202;
assign n_30204 = ~n_30199 & ~n_30203;
assign n_30205 = ~n_30200 & ~n_30204;
assign n_30206 = ~n_30194 & ~n_30198;
assign n_30207 = ~n_30199 & ~n_30206;
assign n_30208 =  x_1870 & ~n_30147;
assign n_30209 = ~n_30195 & ~n_30208;
assign n_30210 = ~n_30193 & ~n_30209;
assign n_30211 = ~n_30194 & ~n_30210;
assign n_30212 = ~n_30149 & ~n_30192;
assign n_30213 = ~n_30193 & ~n_30212;
assign n_30214 =  x_1872 & ~n_30145;
assign n_30215 = ~n_30146 & ~n_30214;
assign n_30216 = ~n_30191 & ~n_30215;
assign n_30217 = ~n_30192 & ~n_30216;
assign n_30218 = ~n_30151 & ~n_30190;
assign n_30219 = ~n_30191 & ~n_30218;
assign n_30220 =  x_1874 & ~n_30143;
assign n_30221 = ~n_30144 & ~n_30220;
assign n_30222 = ~n_30189 & ~n_30221;
assign n_30223 = ~n_30190 & ~n_30222;
assign n_30224 = ~n_30153 & ~n_30188;
assign n_30225 = ~n_30189 & ~n_30224;
assign n_30226 =  x_1876 & ~n_30141;
assign n_30227 = ~n_30142 & ~n_30226;
assign n_30228 = ~n_30187 & ~n_30227;
assign n_30229 = ~n_30188 & ~n_30228;
assign n_30230 = ~n_30155 & ~n_30186;
assign n_30231 = ~n_30187 & ~n_30230;
assign n_30232 =  x_1878 & ~n_30139;
assign n_30233 = ~n_30140 & ~n_30232;
assign n_30234 = ~n_30185 & ~n_30233;
assign n_30235 = ~n_30186 & ~n_30234;
assign n_30236 = ~n_30157 & ~n_30184;
assign n_30237 = ~n_30185 & ~n_30236;
assign n_30238 =  x_1880 & ~n_30137;
assign n_30239 = ~n_30138 & ~n_30238;
assign n_30240 = ~n_30183 & ~n_30239;
assign n_30241 = ~n_30184 & ~n_30240;
assign n_30242 = ~n_30159 & ~n_30182;
assign n_30243 = ~n_30183 & ~n_30242;
assign n_30244 =  x_1882 & ~n_30135;
assign n_30245 = ~n_30136 & ~n_30244;
assign n_30246 = ~n_30181 & ~n_30245;
assign n_30247 = ~n_30182 & ~n_30246;
assign n_30248 = ~n_30161 & ~n_30180;
assign n_30249 = ~n_30181 & ~n_30248;
assign n_30250 =  x_1884 & ~n_30133;
assign n_30251 = ~n_30134 & ~n_30250;
assign n_30252 = ~n_30179 & ~n_30251;
assign n_30253 = ~n_30180 & ~n_30252;
assign n_30254 = ~n_30163 & ~n_30178;
assign n_30255 = ~n_30179 & ~n_30254;
assign n_30256 =  x_1886 & ~n_30131;
assign n_30257 = ~n_30132 & ~n_30256;
assign n_30258 = ~n_30177 & ~n_30257;
assign n_30259 = ~n_30178 & ~n_30258;
assign n_30260 = ~n_30165 & ~n_30176;
assign n_30261 = ~n_30177 & ~n_30260;
assign n_30262 =  x_1888 & ~n_30129;
assign n_30263 = ~n_30130 & ~n_30262;
assign n_30264 = ~n_30175 & ~n_30263;
assign n_30265 = ~n_30176 & ~n_30264;
assign n_30266 = ~n_30167 & ~n_30174;
assign n_30267 = ~n_30175 & ~n_30266;
assign n_30268 =  x_1890 & ~n_30127;
assign n_30269 = ~n_30128 & ~n_30268;
assign n_30270 = ~n_30173 & ~n_30269;
assign n_30271 = ~n_30174 & ~n_30270;
assign n_30272 = ~n_30169 & ~n_30172;
assign n_30273 = ~n_30173 & ~n_30272;
assign n_30274 = ~n_30125 & ~n_30171;
assign n_30275 =  x_1892 & ~n_30274;
assign n_30276 = ~x_1892 &  n_30274;
assign n_30277 = ~n_30275 & ~n_30276;
assign n_30278 =  x_1893 & ~n_30123;
assign n_30279 =  n_30274 & ~n_30278;
assign n_30280 =  x_1895 & ~n_30121;
assign n_30281 = ~n_30122 & ~n_30280;
assign n_30282 = ~x_1865 & ~x_1897;
assign n_30283 =  x_1866 & ~x_1898;
assign n_30284 =  x_1865 &  x_1897;
assign n_30285 = ~n_30283 & ~n_30284;
assign n_30286 = ~n_30282 & ~n_30285;
assign n_30287 = ~x_1864 & ~n_30286;
assign n_30288 =  x_1896 & ~x_1897;
assign n_30289 = ~x_1896 &  x_1897;
assign n_30290 = ~n_30288 & ~n_30289;
assign n_30291 =  x_1864 &  n_30286;
assign n_30292 =  n_30290 & ~n_30291;
assign n_30293 = ~n_30287 & ~n_30292;
assign n_30294 = ~n_30281 & ~n_30293;
assign n_30295 =  n_30281 &  n_30293;
assign n_30296 = ~x_1863 & ~n_30295;
assign n_30297 = ~n_30294 & ~n_30296;
assign n_30298 =  x_1894 & ~n_30122;
assign n_30299 = ~n_30123 & ~n_30298;
assign n_30300 = ~n_30297 & ~n_30299;
assign n_30301 =  n_30297 &  n_30299;
assign n_30302 = ~x_1862 & ~n_30301;
assign n_30303 = ~n_30300 & ~n_30302;
assign n_30304 = ~n_30279 & ~n_30303;
assign n_30305 =  n_30279 &  n_30303;
assign n_30306 = ~x_1861 & ~n_30305;
assign n_30307 = ~n_30304 & ~n_30306;
assign n_30308 =  n_30277 & ~n_30307;
assign n_30309 = ~n_30277 &  n_30307;
assign n_30310 = ~x_1860 & ~n_30309;
assign n_30311 = ~n_30308 & ~n_30310;
assign n_30312 = ~n_30273 & ~n_30311;
assign n_30313 =  n_30273 &  n_30311;
assign n_30314 = ~x_1859 & ~n_30313;
assign n_30315 = ~n_30312 & ~n_30314;
assign n_30316 = ~n_30271 & ~n_30315;
assign n_30317 =  n_30271 &  n_30315;
assign n_30318 = ~x_1858 & ~n_30317;
assign n_30319 = ~n_30316 & ~n_30318;
assign n_30320 = ~n_30267 & ~n_30319;
assign n_30321 =  n_30267 &  n_30319;
assign n_30322 = ~x_1857 & ~n_30321;
assign n_30323 = ~n_30320 & ~n_30322;
assign n_30324 = ~n_30265 & ~n_30323;
assign n_30325 =  n_30265 &  n_30323;
assign n_30326 = ~x_1856 & ~n_30325;
assign n_30327 = ~n_30324 & ~n_30326;
assign n_30328 = ~n_30261 & ~n_30327;
assign n_30329 =  n_30261 &  n_30327;
assign n_30330 = ~x_1855 & ~n_30329;
assign n_30331 = ~n_30328 & ~n_30330;
assign n_30332 = ~n_30259 & ~n_30331;
assign n_30333 =  n_30259 &  n_30331;
assign n_30334 = ~x_1854 & ~n_30333;
assign n_30335 = ~n_30332 & ~n_30334;
assign n_30336 = ~n_30255 & ~n_30335;
assign n_30337 =  n_30255 &  n_30335;
assign n_30338 = ~x_1853 & ~n_30337;
assign n_30339 = ~n_30336 & ~n_30338;
assign n_30340 = ~n_30253 & ~n_30339;
assign n_30341 =  n_30253 &  n_30339;
assign n_30342 = ~x_1852 & ~n_30341;
assign n_30343 = ~n_30340 & ~n_30342;
assign n_30344 = ~n_30249 & ~n_30343;
assign n_30345 =  n_30249 &  n_30343;
assign n_30346 = ~x_1851 & ~n_30345;
assign n_30347 = ~n_30344 & ~n_30346;
assign n_30348 = ~n_30247 & ~n_30347;
assign n_30349 =  n_30247 &  n_30347;
assign n_30350 = ~x_1850 & ~n_30349;
assign n_30351 = ~n_30348 & ~n_30350;
assign n_30352 = ~n_30243 & ~n_30351;
assign n_30353 =  n_30243 &  n_30351;
assign n_30354 = ~x_1849 & ~n_30353;
assign n_30355 = ~n_30352 & ~n_30354;
assign n_30356 = ~n_30241 & ~n_30355;
assign n_30357 =  n_30241 &  n_30355;
assign n_30358 = ~x_1848 & ~n_30357;
assign n_30359 = ~n_30356 & ~n_30358;
assign n_30360 = ~n_30237 & ~n_30359;
assign n_30361 =  n_30237 &  n_30359;
assign n_30362 = ~x_1847 & ~n_30361;
assign n_30363 = ~n_30360 & ~n_30362;
assign n_30364 = ~n_30235 & ~n_30363;
assign n_30365 =  n_30235 &  n_30363;
assign n_30366 = ~x_1846 & ~n_30365;
assign n_30367 = ~n_30364 & ~n_30366;
assign n_30368 = ~n_30231 & ~n_30367;
assign n_30369 =  n_30231 &  n_30367;
assign n_30370 = ~x_1845 & ~n_30369;
assign n_30371 = ~n_30368 & ~n_30370;
assign n_30372 = ~n_30229 & ~n_30371;
assign n_30373 =  n_30229 &  n_30371;
assign n_30374 = ~x_1844 & ~n_30373;
assign n_30375 = ~n_30372 & ~n_30374;
assign n_30376 = ~n_30225 & ~n_30375;
assign n_30377 =  n_30225 &  n_30375;
assign n_30378 = ~x_1843 & ~n_30377;
assign n_30379 = ~n_30376 & ~n_30378;
assign n_30380 = ~n_30223 & ~n_30379;
assign n_30381 =  n_30223 &  n_30379;
assign n_30382 = ~x_1842 & ~n_30381;
assign n_30383 = ~n_30380 & ~n_30382;
assign n_30384 = ~n_30219 & ~n_30383;
assign n_30385 =  n_30219 &  n_30383;
assign n_30386 = ~x_1841 & ~n_30385;
assign n_30387 = ~n_30384 & ~n_30386;
assign n_30388 = ~n_30217 & ~n_30387;
assign n_30389 =  n_30217 &  n_30387;
assign n_30390 = ~x_1840 & ~n_30389;
assign n_30391 = ~n_30388 & ~n_30390;
assign n_30392 = ~n_30213 & ~n_30391;
assign n_30393 =  n_30213 &  n_30391;
assign n_30394 = ~x_1839 & ~n_30393;
assign n_30395 = ~n_30392 & ~n_30394;
assign n_30396 = ~n_30211 & ~n_30395;
assign n_30397 =  n_30211 &  n_30395;
assign n_30398 = ~x_1838 & ~n_30397;
assign n_30399 = ~n_30396 & ~n_30398;
assign n_30400 = ~n_30207 & ~n_30399;
assign n_30401 =  n_30207 &  n_30399;
assign n_30402 = ~x_1837 & ~n_30401;
assign n_30403 = ~n_30400 & ~n_30402;
assign n_30404 =  n_30205 &  n_30403;
assign n_30405 = ~n_30205 & ~n_30403;
assign n_30406 =  x_1836 & ~n_30405;
assign n_30407 =  n_30404 & ~n_30406;
assign n_30408 = ~n_30404 &  n_30406;
assign n_30409 = ~n_30407 & ~n_30408;
assign n_30410 = ~x_1867 & ~n_30201;
assign n_30411 = ~n_30200 &  n_30410;
assign n_30412 = ~x_1835 & ~n_30411;
assign n_30413 =  x_1867 &  n_30201;
assign n_30414 = ~n_30410 & ~n_30413;
assign n_30415 = ~n_30200 &  n_30414;
assign n_30416 =  n_30200 & ~n_30414;
assign n_30417 = ~n_30415 & ~n_30416;
assign n_30418 =  x_1835 &  n_30417;
assign n_30419 = ~n_30412 & ~n_30418;
assign n_30420 = ~n_30409 &  n_30419;
assign n_30421 = ~x_1835 & ~n_30417;
assign n_30422 = ~n_30418 & ~n_30421;
assign n_30423 = ~x_1836 & ~n_30411;
assign n_30424 = ~n_30422 &  n_30423;
assign n_30425 =  n_30405 &  n_30424;
assign n_30426 = ~n_30420 & ~n_30425;
assign n_30427 = ~n_30400 & ~n_30401;
assign n_30428 = ~x_1837 &  n_30427;
assign n_30429 =  x_1837 & ~n_30427;
assign n_30430 = ~n_30396 & ~n_30397;
assign n_30431 =  x_1838 &  n_30430;
assign n_30432 = ~x_1838 & ~n_30430;
assign n_30433 = ~n_30431 & ~n_30432;
assign n_30434 = ~n_30392 & ~n_30393;
assign n_30435 =  x_1839 &  n_30434;
assign n_30436 = ~x_1839 & ~n_30434;
assign n_30437 = ~n_30435 & ~n_30436;
assign n_30438 = ~n_30388 & ~n_30389;
assign n_30439 =  x_1840 &  n_30438;
assign n_30440 = ~x_1840 & ~n_30438;
assign n_30441 = ~n_30439 & ~n_30440;
assign n_30442 = ~n_30384 & ~n_30385;
assign n_30443 =  x_1841 &  n_30442;
assign n_30444 = ~x_1841 & ~n_30442;
assign n_30445 = ~n_30443 & ~n_30444;
assign n_30446 = ~n_30380 & ~n_30381;
assign n_30447 =  x_1842 &  n_30446;
assign n_30448 = ~x_1842 & ~n_30446;
assign n_30449 = ~n_30447 & ~n_30448;
assign n_30450 = ~n_30376 & ~n_30377;
assign n_30451 =  x_1843 &  n_30450;
assign n_30452 = ~x_1843 & ~n_30450;
assign n_30453 = ~n_30451 & ~n_30452;
assign n_30454 = ~n_30372 & ~n_30373;
assign n_30455 =  x_1844 &  n_30454;
assign n_30456 = ~x_1844 & ~n_30454;
assign n_30457 = ~n_30455 & ~n_30456;
assign n_30458 = ~n_30368 & ~n_30369;
assign n_30459 =  x_1845 &  n_30458;
assign n_30460 = ~x_1845 & ~n_30458;
assign n_30461 = ~n_30459 & ~n_30460;
assign n_30462 = ~n_30364 & ~n_30365;
assign n_30463 =  x_1846 &  n_30462;
assign n_30464 = ~x_1846 & ~n_30462;
assign n_30465 = ~n_30463 & ~n_30464;
assign n_30466 = ~n_30360 & ~n_30361;
assign n_30467 =  x_1847 &  n_30466;
assign n_30468 = ~x_1847 & ~n_30466;
assign n_30469 = ~n_30467 & ~n_30468;
assign n_30470 = ~n_30356 & ~n_30357;
assign n_30471 =  x_1848 &  n_30470;
assign n_30472 = ~x_1848 & ~n_30470;
assign n_30473 = ~n_30471 & ~n_30472;
assign n_30474 = ~n_30352 & ~n_30353;
assign n_30475 =  x_1849 &  n_30474;
assign n_30476 = ~x_1849 & ~n_30474;
assign n_30477 = ~n_30475 & ~n_30476;
assign n_30478 = ~n_30348 & ~n_30349;
assign n_30479 =  x_1850 &  n_30478;
assign n_30480 = ~x_1850 & ~n_30478;
assign n_30481 = ~n_30479 & ~n_30480;
assign n_30482 = ~n_30344 & ~n_30345;
assign n_30483 =  x_1851 &  n_30482;
assign n_30484 = ~x_1851 & ~n_30482;
assign n_30485 = ~n_30483 & ~n_30484;
assign n_30486 = ~n_30340 & ~n_30341;
assign n_30487 =  x_1852 &  n_30486;
assign n_30488 = ~x_1852 & ~n_30486;
assign n_30489 = ~n_30487 & ~n_30488;
assign n_30490 = ~n_30336 & ~n_30337;
assign n_30491 =  x_1853 &  n_30490;
assign n_30492 = ~x_1853 & ~n_30490;
assign n_30493 = ~n_30491 & ~n_30492;
assign n_30494 = ~n_30332 & ~n_30333;
assign n_30495 =  x_1854 &  n_30494;
assign n_30496 = ~x_1854 & ~n_30494;
assign n_30497 = ~n_30495 & ~n_30496;
assign n_30498 = ~n_30328 & ~n_30329;
assign n_30499 =  x_1855 &  n_30498;
assign n_30500 = ~x_1855 & ~n_30498;
assign n_30501 = ~n_30499 & ~n_30500;
assign n_30502 = ~n_30324 & ~n_30325;
assign n_30503 =  x_1856 &  n_30502;
assign n_30504 = ~x_1856 & ~n_30502;
assign n_30505 = ~n_30503 & ~n_30504;
assign n_30506 = ~n_30320 & ~n_30321;
assign n_30507 =  x_1857 &  n_30506;
assign n_30508 = ~x_1857 & ~n_30506;
assign n_30509 = ~n_30507 & ~n_30508;
assign n_30510 = ~n_30316 & ~n_30317;
assign n_30511 =  x_1858 &  n_30510;
assign n_30512 = ~x_1858 & ~n_30510;
assign n_30513 = ~n_30511 & ~n_30512;
assign n_30514 = ~n_30312 & ~n_30313;
assign n_30515 =  x_1859 &  n_30514;
assign n_30516 = ~x_1859 & ~n_30514;
assign n_30517 = ~n_30515 & ~n_30516;
assign n_30518 = ~n_30308 & ~n_30309;
assign n_30519 =  x_1860 &  n_30518;
assign n_30520 = ~x_1860 & ~n_30518;
assign n_30521 = ~n_30519 & ~n_30520;
assign n_30522 = ~n_30304 & ~n_30305;
assign n_30523 =  x_1861 &  n_30522;
assign n_30524 = ~x_1861 & ~n_30522;
assign n_30525 = ~n_30523 & ~n_30524;
assign n_30526 = ~n_30300 & ~n_30301;
assign n_30527 =  x_1862 &  n_30526;
assign n_30528 = ~x_1862 & ~n_30526;
assign n_30529 = ~n_30527 & ~n_30528;
assign n_30530 = ~n_30294 & ~n_30295;
assign n_30531 =  x_1863 &  n_30530;
assign n_30532 = ~x_1863 & ~n_30530;
assign n_30533 = ~n_30531 & ~n_30532;
assign n_30534 = ~n_30287 & ~n_30291;
assign n_30535 = ~n_30290 & ~n_30534;
assign n_30536 = ~n_30287 &  n_30292;
assign n_30537 = ~n_30282 & ~n_30284;
assign n_30538 = ~x_1866 &  x_1898;
assign n_30539 = ~n_30283 & ~n_30538;
assign n_30540 = ~n_30537 &  n_30539;
assign n_30541 = ~n_30536 &  n_30540;
assign n_30542 = ~n_30535 &  n_30541;
assign n_30543 = ~n_30533 &  n_30542;
assign n_30544 = ~n_30529 &  n_30543;
assign n_30545 = ~n_30525 &  n_30544;
assign n_30546 = ~n_30521 &  n_30545;
assign n_30547 = ~n_30517 &  n_30546;
assign n_30548 = ~n_30513 &  n_30547;
assign n_30549 = ~n_30509 &  n_30548;
assign n_30550 = ~n_30505 &  n_30549;
assign n_30551 = ~n_30501 &  n_30550;
assign n_30552 = ~n_30497 &  n_30551;
assign n_30553 = ~n_30493 &  n_30552;
assign n_30554 = ~n_30489 &  n_30553;
assign n_30555 = ~n_30485 &  n_30554;
assign n_30556 = ~n_30481 &  n_30555;
assign n_30557 = ~n_30477 &  n_30556;
assign n_30558 = ~n_30473 &  n_30557;
assign n_30559 = ~n_30469 &  n_30558;
assign n_30560 = ~n_30465 &  n_30559;
assign n_30561 = ~n_30461 &  n_30560;
assign n_30562 = ~n_30457 &  n_30561;
assign n_30563 = ~n_30453 &  n_30562;
assign n_30564 = ~n_30449 &  n_30563;
assign n_30565 = ~n_30445 &  n_30564;
assign n_30566 = ~n_30441 &  n_30565;
assign n_30567 = ~n_30437 &  n_30566;
assign n_30568 = ~n_30433 &  n_30567;
assign n_30569 = ~n_30429 &  n_30568;
assign n_30570 = ~n_30428 &  n_30569;
assign n_30571 = ~n_30426 &  n_30570;
assign n_30572 =  n_25775 & ~n_30571;
assign n_30573 =  n_8818 &  n_28634;
assign n_30574 = ~n_29440 & ~n_27405;
assign n_30575 = ~n_30573 &  n_30574;
assign n_30576 = ~n_28571 & ~n_28635;
assign n_30577 =  n_30575 &  n_30576;
assign n_30578 =  n_29248 &  n_28588;
assign n_30579 =  n_30577 &  n_30578;
assign n_30580 = ~n_27264 &  n_29659;
assign n_30581 = ~n_27412 &  n_30580;
assign n_30582 = ~n_28617 &  n_28601;
assign n_30583 =  n_8060 &  n_29255;
assign n_30584 =  n_27976 &  n_30583;
assign n_30585 = ~n_30584 & ~n_29078;
assign n_30586 = ~n_28648 & ~n_27933;
assign n_30587 =  n_30585 &  n_30586;
assign n_30588 =  n_28938 &  n_30587;
assign n_30589 = ~n_29491 &  n_29327;
assign n_30590 =  n_28537 &  n_28029;
assign n_30591 = ~n_30590 &  n_28646;
assign n_30592 =  n_30589 &  n_30591;
assign n_30593 =  n_30588 &  n_30592;
assign n_30594 = ~n_28942 & ~n_28653;
assign n_30595 =  n_30594 &  n_28643;
assign n_30596 =  n_30593 &  n_30595;
assign n_30597 = ~n_24802 & ~n_28742;
assign n_30598 =  n_30597 &  n_29339;
assign n_30599 =  n_30598 &  n_28954;
assign n_30600 =  n_29639 &  n_30599;
assign n_30601 =  n_29347 &  n_29649;
assign n_30602 =  n_30600 &  n_30601;
assign n_30603 = ~n_29298 & ~n_28013;
assign n_30604 =  n_27259 &  n_1906;
assign n_30605 = ~n_30604 & ~n_6529;
assign n_30606 = ~n_29380 & ~n_4058;
assign n_30607 =  n_6527 &  n_6533;
assign n_30608 = ~n_30607 & ~n_3863;
assign n_30609 =  n_30606 &  n_30608;
assign n_30610 =  n_30605 &  n_30609;
assign n_30611 =  n_30603 &  n_30610;
assign n_30612 =  x_37 &  n_29230;
assign n_30613 = ~n_29097 & ~n_30612;
assign n_30614 = ~n_28752 &  n_30613;
assign n_30615 = ~n_24607 & ~n_16334;
assign n_30616 =  n_27424 &  n_186;
assign n_30617 = ~n_30616 & ~n_16528;
assign n_30618 =  n_30615 &  n_30617;
assign n_30619 =  n_30614 &  n_30618;
assign n_30620 =  n_29199 & ~n_28911;
assign n_30621 =  n_30619 &  n_30620;
assign n_30622 =  n_30611 &  n_30621;
assign n_30623 = ~n_28865 & ~n_27909;
assign n_30624 = ~n_27584 &  n_30623;
assign n_30625 =  n_28871 &  n_29617;
assign n_30626 =  n_30624 &  n_30625;
assign n_30627 =  n_28740 &  n_29165;
assign n_30628 = ~n_28999 & ~n_29014;
assign n_30629 = ~n_28238 &  n_30628;
assign n_30630 = ~n_2304 &  n_29516;
assign n_30631 =  n_30629 &  n_30630;
assign n_30632 =  n_30627 &  n_30631;
assign n_30633 =  n_30626 &  n_30632;
assign n_30634 =  n_30622 &  n_30633;
assign n_30635 =  n_28436 &  n_28820;
assign n_30636 = ~n_28832 & ~n_30635;
assign n_30637 = ~n_28688 & ~n_28866;
assign n_30638 =  n_30636 &  n_30637;
assign n_30639 = ~n_28930 & ~n_28782;
assign n_30640 =  x_38 &  n_24801;
assign n_30641 =  n_785 &  n_30640;
assign n_30642 = ~n_30641 & ~n_28692;
assign n_30643 =  n_30642 &  n_29354;
assign n_30644 =  n_30639 &  n_30643;
assign n_30645 =  n_30638 &  n_30644;
assign n_30646 = ~n_28788 & ~n_19946;
assign n_30647 =  n_28428 &  n_30646;
assign n_30648 = ~n_29411 &  n_30647;
assign n_30649 = ~x_735 & ~x_736;
assign n_30650 = ~x_737 & ~x_738;
assign n_30651 =  n_30649 &  n_30650;
assign n_30652 = ~x_731 & ~x_732;
assign n_30653 = ~x_733 & ~x_734;
assign n_30654 =  n_30652 &  n_30653;
assign n_30655 =  n_30651 &  n_30654;
assign n_30656 = ~x_743 & ~x_744;
assign n_30657 = ~x_745 & ~x_746;
assign n_30658 =  n_30656 &  n_30657;
assign n_30659 = ~x_739 & ~x_740;
assign n_30660 = ~x_741 & ~x_742;
assign n_30661 =  n_30659 &  n_30660;
assign n_30662 =  n_30658 &  n_30661;
assign n_30663 =  n_30655 &  n_30662;
assign n_30664 = ~x_719 & ~x_720;
assign n_30665 = ~x_721 & ~x_722;
assign n_30666 =  n_30664 &  n_30665;
assign n_30667 = ~x_715 & ~x_716;
assign n_30668 = ~x_717 & ~x_718;
assign n_30669 =  n_30667 &  n_30668;
assign n_30670 =  n_30666 &  n_30669;
assign n_30671 = ~x_727 & ~x_728;
assign n_30672 = ~x_729 & ~x_730;
assign n_30673 =  n_30671 &  n_30672;
assign n_30674 = ~x_723 & ~x_724;
assign n_30675 = ~x_725 & ~x_726;
assign n_30676 =  n_30674 &  n_30675;
assign n_30677 =  n_30673 &  n_30676;
assign n_30678 =  n_30670 &  n_30677;
assign n_30679 =  n_30663 &  n_30678;
assign n_30680 =  n_28829 &  n_30679;
assign n_30681 = ~n_30680 & ~n_28166;
assign n_30682 =  n_29190 &  n_28835;
assign n_30683 =  n_30681 &  n_30682;
assign n_30684 =  n_30648 &  n_30683;
assign n_30685 =  n_30645 &  n_30684;
assign n_30686 = ~n_28461 & ~n_28728;
assign n_30687 = ~n_29307 & ~n_5197;
assign n_30688 =  n_30686 &  n_30687;
assign n_30689 = ~n_28722 & ~n_20139;
assign n_30690 = ~n_27550 &  n_30689;
assign n_30691 = ~n_29486 & ~n_28915;
assign n_30692 =  n_30690 &  n_30691;
assign n_30693 =  n_30688 &  n_30692;
assign n_30694 = ~n_20332 & ~n_27934;
assign n_30695 = ~n_28780 & ~n_28828;
assign n_30696 =  n_30694 &  n_30695;
assign n_30697 = ~n_22538 & ~n_391;
assign n_30698 = ~n_28326 & ~n_5192;
assign n_30699 =  n_30697 &  n_30698;
assign n_30700 =  n_30696 &  n_30699;
assign n_30701 =  n_30693 &  n_30700;
assign n_30702 = ~n_25776 & ~n_18446;
assign n_30703 = ~n_28219 &  n_30702;
assign n_30704 =  n_28980 & ~n_28736;
assign n_30705 =  n_30703 &  n_30704;
assign n_30706 = ~n_28589 & ~n_28471;
assign n_30707 =  n_29110 &  n_30706;
assign n_30708 = ~n_28451 & ~n_29505;
assign n_30709 =  n_30708 & ~n_28773;
assign n_30710 =  n_30707 &  n_30709;
assign n_30711 =  n_30705 &  n_30710;
assign n_30712 =  n_30701 &  n_30711;
assign n_30713 =  n_30685 &  n_30712;
assign n_30714 =  n_30634 &  n_30713;
assign n_30715 = ~n_28447 & ~n_29396;
assign n_30716 = ~n_28694 & ~n_28523;
assign n_30717 = ~n_29622 &  n_30716;
assign n_30718 =  n_30715 &  n_30717;
assign n_30719 =  n_27818 &  n_30718;
assign n_30720 =  n_27605 &  n_29333;
assign n_30721 =  n_30719 &  n_30720;
assign n_30722 = ~n_28872 &  n_29609;
assign n_30723 =  n_28427 &  n_29612;
assign n_30724 =  n_30722 &  n_30723;
assign n_30725 =  n_27979 &  n_30724;
assign n_30726 = ~n_28924 & ~n_28926;
assign n_30727 =  n_30725 &  n_30726;
assign n_30728 =  n_30721 &  n_30727;
assign n_30729 =  n_30714 &  n_30728;
assign n_30730 =  n_30602 &  n_30729;
assign n_30731 =  n_30596 &  n_30730;
assign n_30732 = ~n_27426 &  n_30731;
assign n_30733 = ~n_27254 &  n_28525;
assign n_30734 = ~n_27418 & ~n_30733;
assign n_30735 =  n_30732 &  n_30734;
assign n_30736 =  n_30582 &  n_30735;
assign n_30737 =  n_30581 &  n_30736;
assign n_30738 =  n_29485 &  n_30737;
assign n_30739 =  n_30579 &  n_30738;
assign n_30740 = ~n_30572 &  n_30739;
assign n_30741 = ~n_30120 &  n_30740;
assign n_30742 =  x_37 & ~n_30741;
assign n_30743 = ~x_37 &  n_30741;
assign n_30744 = ~n_30742 & ~n_30743;
assign n_30745 =  n_28550 & ~n_30119;
assign n_30746 = ~n_29638 & ~n_27749;
assign n_30747 =  n_28995 &  n_29605;
assign n_30748 =  n_30746 &  n_30747;
assign n_30749 =  n_28329 &  n_30623;
assign n_30750 = ~n_28026 &  n_29615;
assign n_30751 =  n_30749 &  n_30750;
assign n_30752 =  n_28779 &  n_29176;
assign n_30753 = ~n_28341 &  n_29302;
assign n_30754 =  n_30752 &  n_30753;
assign n_30755 =  n_30751 &  n_30754;
assign n_30756 = ~n_1907 & ~n_2102;
assign n_30757 = ~n_22266 &  n_30756;
assign n_30758 =  n_29110 &  n_30757;
assign n_30759 =  n_28548 &  n_30758;
assign n_30760 =  n_28312 & ~n_28040;
assign n_30761 =  n_29304 &  n_30760;
assign n_30762 =  n_30759 &  n_30761;
assign n_30763 =  n_30755 &  n_30762;
assign n_30764 =  n_30748 &  n_30763;
assign n_30765 =  n_30718 &  n_28858;
assign n_30766 =  n_29264 &  n_27591;
assign n_30767 =  n_30765 &  n_30766;
assign n_30768 =  n_28860 &  n_27827;
assign n_30769 =  n_28975 &  n_29299;
assign n_30770 =  n_30768 &  n_30769;
assign n_30771 =  n_30767 &  n_30770;
assign n_30772 =  n_30764 &  n_30771;
assign n_30773 =  n_29057 &  n_29592;
assign n_30774 = ~n_29324 &  n_28785;
assign n_30775 =  n_30773 &  n_30774;
assign n_30776 = ~n_27834 &  n_30775;
assign n_30777 = ~n_29080 & ~n_28243;
assign n_30778 = ~n_29646 &  n_30777;
assign n_30779 = ~n_28846 &  n_30778;
assign n_30780 =  n_30779 &  n_29342;
assign n_30781 =  n_30776 &  n_30780;
assign n_30782 = ~n_29353 & ~n_28697;
assign n_30783 = ~n_1707 & ~n_24801;
assign n_30784 =  n_191 & ~n_30783;
assign n_30785 = ~n_28126 & ~n_27670;
assign n_30786 = ~n_30784 &  n_30785;
assign n_30787 =  n_30782 &  n_30786;
assign n_30788 =  n_28212 & ~n_28986;
assign n_30789 =  n_30787 &  n_30788;
assign n_30790 = ~n_29101 & ~n_29419;
assign n_30791 = ~n_3863 & ~n_6534;
assign n_30792 =  n_30790 &  n_30791;
assign n_30793 = ~n_29200 & ~n_21879;
assign n_30794 = ~n_28914 & ~n_4252;
assign n_30795 =  n_30793 &  n_30794;
assign n_30796 =  n_30792 &  n_30795;
assign n_30797 =  n_30789 &  n_30796;
assign n_30798 = ~n_391 & ~n_786;
assign n_30799 = ~n_29626 &  n_30798;
assign n_30800 = ~n_27912 & ~n_29009;
assign n_30801 =  n_30799 &  n_30800;
assign n_30802 = ~n_28771 & ~n_28529;
assign n_30803 =  n_28565 &  n_1315;
assign n_30804 =  n_30606 & ~n_30803;
assign n_30805 =  n_30802 &  n_30804;
assign n_30806 =  n_30801 &  n_30805;
assign n_30807 =  n_30797 &  n_30806;
assign n_30808 =  n_29251 &  n_29422;
assign n_30809 = ~n_29623 & ~n_27916;
assign n_30810 = ~n_18434 &  n_30809;
assign n_30811 =  n_28848 &  n_30810;
assign n_30812 =  n_30808 &  n_30811;
assign n_30813 = ~n_13021 & ~n_25776;
assign n_30814 = ~n_2304 & ~n_27708;
assign n_30815 =  n_30813 &  n_30814;
assign n_30816 = ~n_28453 & ~n_6531;
assign n_30817 = ~n_28114 & ~n_18440;
assign n_30818 =  n_30816 &  n_30817;
assign n_30819 =  n_30815 &  n_30818;
assign n_30820 =  n_1 &  n_13015;
assign n_30821 =  n_28751 & ~n_30820;
assign n_30822 = ~n_20914 &  n_30821;
assign n_30823 = ~n_29188 & ~n_28027;
assign n_30824 =  n_29389 &  n_28539;
assign n_30825 =  n_30823 &  n_30824;
assign n_30826 =  n_30822 &  n_30825;
assign n_30827 =  n_30819 &  n_30826;
assign n_30828 =  n_30812 &  n_30827;
assign n_30829 =  n_30807 &  n_30828;
assign n_30830 =  n_29075 &  n_28513;
assign n_30831 = ~n_29311 &  n_30830;
assign n_30832 =  n_30597 &  n_30831;
assign n_30833 = ~n_29553 & ~n_28947;
assign n_30834 =  n_28737 &  n_30833;
assign n_30835 =  n_28222 &  n_30834;
assign n_30836 =  n_30832 &  n_30835;
assign n_30837 =  n_29086 &  n_30642;
assign n_30838 =  n_29351 & ~n_27841;
assign n_30839 =  n_30837 &  n_30838;
assign n_30840 =  n_29357 &  n_28472;
assign n_30841 = ~n_585 & ~n_1;
assign n_30842 =  n_23892 &  n_30841;
assign n_30843 =  n_29058 & ~n_30842;
assign n_30844 =  n_30840 &  n_30843;
assign n_30845 =  n_30839 &  n_30844;
assign n_30846 = ~n_27933 & ~n_28940;
assign n_30847 =  n_30845 &  n_30846;
assign n_30848 =  n_30836 &  n_30847;
assign n_30849 =  n_30829 &  n_30848;
assign n_30850 =  n_30781 &  n_30849;
assign n_30851 =  n_30772 &  n_30850;
assign n_30852 = ~n_28581 &  n_30851;
assign n_30853 = ~n_28632 & ~n_28587;
assign n_30854 = ~n_28590 &  n_30853;
assign n_30855 =  n_30852 &  n_30854;
assign n_30856 =  n_29218 &  n_29480;
assign n_30857 =  n_30855 &  n_30856;
assign n_30858 =  n_29467 &  n_30857;
assign n_30859 = ~n_29246 &  n_29659;
assign n_30860 = ~n_27254 &  n_28566;
assign n_30861 = ~n_30860 & ~n_28584;
assign n_30862 =  n_28616 &  n_30861;
assign n_30863 =  n_30859 &  n_30862;
assign n_30864 =  n_29446 &  n_28619;
assign n_30865 =  n_30576 &  n_29245;
assign n_30866 =  n_30864 &  n_30865;
assign n_30867 =  n_30863 &  n_30866;
assign n_30868 =  n_30858 &  n_30867;
assign n_30869 = ~n_27129 &  n_30868;
assign n_30870 = ~n_28630 &  n_30869;
assign n_30871 = ~n_30745 &  n_30870;
assign n_30872 =  x_36 & ~n_30871;
assign n_30873 = ~x_36 &  n_30871;
assign n_30874 = ~n_30872 & ~n_30873;
assign n_30875 =  n_28852 &  n_29631;
assign n_30876 =  n_29600 &  n_30875;
assign n_30877 =  n_29603 &  n_30630;
assign n_30878 =  n_30629 &  n_30877;
assign n_30879 =  n_28979 &  n_30810;
assign n_30880 =  n_28981 &  n_28339;
assign n_30881 =  n_30879 &  n_30880;
assign n_30882 =  n_30878 &  n_30881;
assign n_30883 = ~n_28236 &  n_29258;
assign n_30884 =  n_30882 &  n_30883;
assign n_30885 =  n_30876 &  n_30884;
assign n_30886 =  n_30594 &  n_27837;
assign n_30887 =  n_30885 &  n_30886;
assign n_30888 =  n_28784 &  n_29177;
assign n_30889 =  n_29019 &  n_30888;
assign n_30890 = ~n_28024 &  n_30889;
assign n_30891 =  n_29322 &  n_30779;
assign n_30892 =  n_30890 &  n_30891;
assign n_30893 = ~n_29622 & ~n_29070;
assign n_30894 = ~n_26229 &  n_28718;
assign n_30895 =  n_30893 &  n_30894;
assign n_30896 = ~n_15948 & ~n_29101;
assign n_30897 =  n_30896 & ~n_28602;
assign n_30898 = ~n_29396 &  n_28117;
assign n_30899 =  n_30897 &  n_30898;
assign n_30900 =  n_30895 &  n_30899;
assign n_30901 = ~n_27839 & ~n_15755;
assign n_30902 = ~n_28855 &  n_30901;
assign n_30903 =  n_30702 &  n_28830;
assign n_30904 =  n_29073 & ~n_28865;
assign n_30905 =  n_30903 &  n_30904;
assign n_30906 =  n_30902 &  n_30905;
assign n_30907 =  n_30900 &  n_30906;
assign n_30908 =  n_28213 &  n_29010;
assign n_30909 = ~n_29260 &  n_29013;
assign n_30910 =  n_30908 &  n_30909;
assign n_30911 = ~n_9 & ~n_12033;
assign n_30912 = ~n_27934 & ~n_28330;
assign n_30913 =  n_30911 &  n_30912;
assign n_30914 = ~n_4058 & ~n_1317;
assign n_30915 = ~n_8061 &  n_30914;
assign n_30916 = ~n_28451 & ~n_28770;
assign n_30917 =  n_30915 &  n_30916;
assign n_30918 =  n_30913 &  n_30917;
assign n_30919 = ~n_28350 & ~n_984;
assign n_30920 = ~n_28685 & ~n_27840;
assign n_30921 =  n_30919 &  n_30920;
assign n_30922 = ~n_28013 &  n_30921;
assign n_30923 =  n_30918 &  n_30922;
assign n_30924 =  n_30910 &  n_30923;
assign n_30925 =  n_30907 &  n_30924;
assign n_30926 =  n_29168 &  n_30834;
assign n_30927 =  n_30926 &  n_30832;
assign n_30928 =  n_24801 &  n_29297;
assign n_30929 = ~n_29328 & ~n_28948;
assign n_30930 = ~n_30928 &  n_30929;
assign n_30931 = ~n_30584 &  n_30930;
assign n_30932 =  n_29253 &  n_29429;
assign n_30933 =  n_30931 &  n_30932;
assign n_30934 =  n_30927 &  n_30933;
assign n_30935 =  n_30925 &  n_30934;
assign n_30936 =  n_30892 &  n_30935;
assign n_30937 =  n_28934 &  n_30936;
assign n_30938 =  n_30887 &  n_30937;
assign n_30939 = ~n_28572 &  n_30938;
assign n_30940 = ~n_28587 & ~n_29211;
assign n_30941 =  n_30939 &  n_30940;
assign n_30942 = ~n_28618 &  n_27409;
assign n_30943 =  n_30941 &  n_30942;
assign n_30944 =  n_29480 &  n_30859;
assign n_30945 =  n_30943 &  n_30944;
assign n_30946 =  n_29461 &  n_30945;
assign n_30947 =  x_35 & ~n_30946;
assign n_30948 = ~x_35 &  n_30946;
assign n_30949 = ~n_30947 & ~n_30948;
assign n_30950 =  n_29114 &  n_28445;
assign n_30951 =  n_29115 & ~n_23504;
assign n_30952 =  n_30950 &  n_30951;
assign n_30953 =  n_30648 &  n_30952;
assign n_30954 =  n_29202 &  n_30953;
assign n_30955 = ~n_29261 & ~n_23698;
assign n_30956 = ~n_28701 &  n_30955;
assign n_30957 =  n_12420 &  n_27266;
assign n_30958 = ~n_29401 & ~n_30957;
assign n_30959 = ~n_192 & ~n_29219;
assign n_30960 =  n_30958 &  n_30959;
assign n_30961 = ~n_29112 &  n_30960;
assign n_30962 =  n_30782 &  n_30706;
assign n_30963 =  n_30961 &  n_30962;
assign n_30964 =  n_30956 &  n_30963;
assign n_30965 =  n_30759 &  n_30964;
assign n_30966 =  n_28919 &  n_30965;
assign n_30967 =  n_30954 &  n_30966;
assign n_30968 = ~n_28581 &  n_30967;
assign n_30969 = ~n_27426 &  n_30968;
assign n_30970 = ~n_29465 &  n_30969;
assign n_30971 =  n_29218 &  n_30582;
assign n_30972 =  n_30970 &  n_30971;
assign n_30973 =  n_27272 &  n_30972;
assign n_30974 =  n_29488 &  n_30973;
assign n_30975 =  x_33 & ~n_30974;
assign n_30976 = ~x_33 &  n_30974;
assign n_30977 = ~n_30975 & ~n_30976;
assign n_30978 =  n_30715 &  n_29308;
assign n_30979 =  n_28337 &  n_30978;
assign n_30980 =  n_30605 &  n_29558;
assign n_30981 =  n_29561 &  n_30609;
assign n_30982 =  n_30980 &  n_30981;
assign n_30983 =  n_30979 &  n_30982;
assign n_30984 =  n_29254 &  n_29629;
assign n_30985 =  n_30983 &  n_30984;
assign n_30986 =  n_28729 &  n_30708;
assign n_30987 =  n_29394 &  n_30798;
assign n_30988 =  n_30986 &  n_30987;
assign n_30989 =  n_29519 & ~n_28586;
assign n_30990 = ~n_30803 & ~n_29427;
assign n_30991 =  n_30989 &  n_30990;
assign n_30992 =  n_30988 &  n_30991;
assign n_30993 = ~n_28940 &  n_28216;
assign n_30994 =  n_30992 &  n_30993;
assign n_30995 =  n_28988 &  n_28527;
assign n_30996 = ~n_29298 &  n_28990;
assign n_30997 =  n_30995 &  n_30996;
assign n_30998 = ~n_3470 & ~n_25775;
assign n_30999 =  n_30896 &  n_30998;
assign n_31000 = ~n_28602 &  n_28721;
assign n_31001 =  n_30999 &  n_31000;
assign n_31002 = ~n_30641 & ~n_29616;
assign n_31003 = ~n_27592 &  n_31002;
assign n_31004 = ~n_28717 & ~n_28692;
assign n_31005 = ~n_3082 & ~n_27601;
assign n_31006 =  n_31004 &  n_31005;
assign n_31007 =  n_31003 &  n_31006;
assign n_31008 =  n_31001 &  n_31007;
assign n_31009 =  n_30997 &  n_31008;
assign n_31010 =  n_30994 &  n_31009;
assign n_31011 =  n_30985 &  n_31010;
assign n_31012 =  n_30588 &  n_31011;
assign n_31013 =  n_28222 &  n_29164;
assign n_31014 =  n_28118 &  n_28769;
assign n_31015 =  n_31013 &  n_31014;
assign n_31016 =  n_30930 &  n_28776;
assign n_31017 =  n_31016 &  n_29425;
assign n_31018 =  n_31015 &  n_31017;
assign n_31019 =  n_28021 &  n_29065;
assign n_31020 =  n_31018 &  n_31019;
assign n_31021 =  n_29644 &  n_31020;
assign n_31022 =  n_31012 &  n_31021;
assign n_31023 = ~n_28632 &  n_31022;
assign n_31024 =  n_28573 &  n_31023;
assign n_31025 = ~n_29459 &  n_31024;
assign n_31026 =  n_30575 &  n_31025;
assign n_31027 =  n_30863 &  n_31026;
assign n_31028 =  n_29484 &  n_31027;
assign n_31029 = ~n_27129 &  n_31028;
assign n_31030 =  x_34 & ~n_31029;
assign n_31031 = ~x_34 &  n_31029;
assign n_31032 = ~n_31030 & ~n_31031;
assign n_31033 = ~n_30977 & ~n_31032;
assign n_31034 = ~n_30949 &  n_31033;
assign n_31035 = ~n_30874 &  n_31034;
assign n_31036 = ~n_30744 &  n_31035;
assign n_31037 = ~n_29667 &  n_31036;
assign n_31038 = ~n_29479 &  n_31037;
assign n_31039 = ~n_29241 &  n_31038;
assign n_31040 = ~n_28974 &  n_31039;
assign n_31041 = ~n_28629 &  n_31040;
assign n_31042 = ~n_25319 &  n_31041;
assign n_31043 = ~n_25313 &  n_31042;
assign n_31044 = ~n_25307 &  n_31043;
assign n_31045 = ~n_25301 &  n_31044;
assign n_31046 = ~n_25295 &  n_31045;
assign n_31047 = ~n_25289 &  n_31046;
assign n_31048 = ~n_25283 &  n_31047;
assign n_31049 = ~n_25277 &  n_31048;
assign n_31050 = ~n_25271 &  n_31049;
assign n_31051 = ~n_25265 &  n_31050;
assign n_31052 = ~n_25259 &  n_31051;
assign n_31053 = ~n_25253 &  n_31052;
assign n_31054 = ~n_25247 &  n_31053;
assign n_31055 = ~n_25241 &  n_31054;
assign n_31056 = ~n_25235 &  n_31055;
assign n_31057 = ~n_25229 &  n_31056;
assign n_31058 = ~n_25223 &  n_31057;
assign n_31059 = ~n_25217 &  n_31058;
assign n_31060 = ~n_25211 &  n_31059;
assign n_31061 = ~n_25205 &  n_31060;
assign n_31062 = ~n_25199 &  n_31061;
assign n_31063 = ~n_25193 &  n_31062;
assign n_31064 = ~n_25187 &  n_31063;
assign n_31065 = ~n_25181 &  n_31064;
assign n_31066 = ~n_25175 &  n_31065;
assign n_31067 = ~n_25169 &  n_31066;
assign n_31068 = ~n_25163 &  n_31067;
assign n_31069 = ~n_25157 &  n_31068;
assign n_31070 = ~n_25151 &  n_31069;
assign n_31071 = ~n_25145 &  n_31070;
assign n_31072 = ~n_25139 &  n_31071;
assign n_31073 = ~n_25133 &  n_31072;
assign n_31074 = ~n_25127 &  n_31073;
assign n_31075 = ~n_25121 &  n_31074;
assign n_31076 = ~n_25115 &  n_31075;
assign n_31077 = ~n_25109 &  n_31076;
assign n_31078 = ~n_25103 &  n_31077;
assign n_31079 = ~n_25097 &  n_31078;
assign n_31080 = ~n_25091 &  n_31079;
assign n_31081 = ~n_25085 &  n_31080;
assign n_31082 = ~n_25079 &  n_31081;
assign n_31083 = ~n_25073 &  n_31082;
assign n_31084 = ~n_25067 &  n_31083;
assign n_31085 = ~n_25061 &  n_31084;
assign n_31086 = ~n_25055 &  n_31085;
assign n_31087 = ~n_25049 &  n_31086;
assign n_31088 = ~n_25043 &  n_31087;
assign n_31089 = ~n_25037 &  n_31088;
assign n_31090 = ~n_25031 &  n_31089;
assign n_31091 = ~n_25025 &  n_31090;
assign n_31092 = ~n_25019 &  n_31091;
assign n_31093 = ~n_25013 &  n_31092;
assign n_31094 = ~n_25007 &  n_31093;
assign n_31095 = ~n_25001 &  n_31094;
assign n_31096 = ~n_24994 &  n_31095;
assign n_31097 = ~n_24988 &  n_31096;
assign n_31098 = ~n_24982 &  n_31097;
assign n_31099 = ~n_24976 &  n_31098;
assign n_31100 = ~n_24970 &  n_31099;
assign n_31101 = ~n_24964 &  n_31100;
assign n_31102 = ~n_24958 &  n_31101;
assign n_31103 = ~n_24952 &  n_31102;
assign n_31104 = ~n_24946 &  n_31103;
assign n_31105 = ~n_24940 &  n_31104;
assign n_31106 = ~n_24934 &  n_31105;
assign n_31107 = ~n_24928 &  n_31106;
assign n_31108 = ~n_24922 &  n_31107;
assign n_31109 = ~n_24916 &  n_31108;
assign n_31110 = ~n_24910 &  n_31109;
assign n_31111 = ~n_24904 &  n_31110;
assign n_31112 = ~n_24898 &  n_31111;
assign n_31113 = ~n_24892 &  n_31112;
assign n_31114 = ~n_24886 &  n_31113;
assign n_31115 = ~n_24880 &  n_31114;
assign n_31116 = ~n_24874 &  n_31115;
assign n_31117 = ~n_24868 &  n_31116;
assign n_31118 = ~n_24862 &  n_31117;
assign n_31119 = ~n_24856 &  n_31118;
assign n_31120 = ~n_24850 &  n_31119;
assign n_31121 = ~n_24844 &  n_31120;
assign n_31122 = ~n_24838 &  n_31121;
assign n_31123 = ~n_24832 &  n_31122;
assign n_31124 = ~n_24826 &  n_31123;
assign n_31125 = ~n_24820 &  n_31124;
assign n_31126 = ~n_24814 &  n_31125;
assign n_31127 = ~n_24808 &  n_31126;
assign n_31128 = ~n_24800 &  n_31127;
assign n_31129 = ~n_24794 &  n_31128;
assign n_31130 = ~n_24788 &  n_31129;
assign n_31131 = ~n_24782 &  n_31130;
assign n_31132 = ~n_24776 &  n_31131;
assign n_31133 = ~n_24770 &  n_31132;
assign n_31134 = ~n_24764 &  n_31133;
assign n_31135 = ~n_24758 &  n_31134;
assign n_31136 = ~n_24752 &  n_31135;
assign n_31137 = ~n_24746 &  n_31136;
assign n_31138 = ~n_24740 &  n_31137;
assign n_31139 = ~n_24734 &  n_31138;
assign n_31140 = ~n_24728 &  n_31139;
assign n_31141 = ~n_24722 &  n_31140;
assign n_31142 = ~n_24716 &  n_31141;
assign n_31143 = ~n_24710 &  n_31142;
assign n_31144 = ~n_24704 &  n_31143;
assign n_31145 = ~n_24698 &  n_31144;
assign n_31146 = ~n_24692 &  n_31145;
assign n_31147 = ~n_24686 &  n_31146;
assign n_31148 = ~n_24680 &  n_31147;
assign n_31149 = ~n_24674 &  n_31148;
assign n_31150 = ~n_24668 &  n_31149;
assign n_31151 = ~n_24662 &  n_31150;
assign n_31152 = ~n_24656 &  n_31151;
assign n_31153 = ~n_24650 &  n_31152;
assign n_31154 = ~n_24644 &  n_31153;
assign n_31155 = ~n_24638 &  n_31154;
assign n_31156 = ~n_24632 &  n_31155;
assign n_31157 = ~n_24626 &  n_31156;
assign n_31158 = ~n_24620 &  n_31157;
assign n_31159 = ~n_24614 &  n_31158;
assign n_31160 = ~n_24606 &  n_31159;
assign n_31161 = ~n_24600 &  n_31160;
assign n_31162 = ~n_24594 &  n_31161;
assign n_31163 = ~n_24588 &  n_31162;
assign n_31164 = ~n_24582 &  n_31163;
assign n_31165 = ~n_24576 &  n_31164;
assign n_31166 = ~n_24570 &  n_31165;
assign n_31167 = ~n_24564 &  n_31166;
assign n_31168 = ~n_24558 &  n_31167;
assign n_31169 = ~n_24552 &  n_31168;
assign n_31170 = ~n_24546 &  n_31169;
assign n_31171 = ~n_24540 &  n_31170;
assign n_31172 = ~n_24534 &  n_31171;
assign n_31173 = ~n_24528 &  n_31172;
assign n_31174 = ~n_24522 &  n_31173;
assign n_31175 = ~n_24516 &  n_31174;
assign n_31176 = ~n_24510 &  n_31175;
assign n_31177 = ~n_24504 &  n_31176;
assign n_31178 = ~n_24498 &  n_31177;
assign n_31179 = ~n_24492 &  n_31178;
assign n_31180 = ~n_24486 &  n_31179;
assign n_31181 = ~n_24480 &  n_31180;
assign n_31182 = ~n_24474 &  n_31181;
assign n_31183 = ~n_24468 &  n_31182;
assign n_31184 = ~n_24462 &  n_31183;
assign n_31185 = ~n_24456 &  n_31184;
assign n_31186 = ~n_24450 &  n_31185;
assign n_31187 = ~n_24444 &  n_31186;
assign n_31188 = ~n_24438 &  n_31187;
assign n_31189 = ~n_24432 &  n_31188;
assign n_31190 = ~n_24426 &  n_31189;
assign n_31191 = ~n_24420 &  n_31190;
assign n_31192 = ~n_24412 &  n_31191;
assign n_31193 = ~n_24406 &  n_31192;
assign n_31194 = ~n_24400 &  n_31193;
assign n_31195 = ~n_24394 &  n_31194;
assign n_31196 = ~n_24388 &  n_31195;
assign n_31197 = ~n_24382 &  n_31196;
assign n_31198 = ~n_24376 &  n_31197;
assign n_31199 = ~n_24370 &  n_31198;
assign n_31200 = ~n_24364 &  n_31199;
assign n_31201 = ~n_24358 &  n_31200;
assign n_31202 = ~n_24352 &  n_31201;
assign n_31203 = ~n_24346 &  n_31202;
assign n_31204 = ~n_24340 &  n_31203;
assign n_31205 = ~n_24334 &  n_31204;
assign n_31206 = ~n_24328 &  n_31205;
assign n_31207 = ~n_24322 &  n_31206;
assign n_31208 = ~n_24316 &  n_31207;
assign n_31209 = ~n_24310 &  n_31208;
assign n_31210 = ~n_24304 &  n_31209;
assign n_31211 = ~n_24298 &  n_31210;
assign n_31212 = ~n_24292 &  n_31211;
assign n_31213 = ~n_24286 &  n_31212;
assign n_31214 = ~n_24280 &  n_31213;
assign n_31215 = ~n_24274 &  n_31214;
assign n_31216 = ~n_24268 &  n_31215;
assign n_31217 = ~n_24262 &  n_31216;
assign n_31218 = ~n_24256 &  n_31217;
assign n_31219 = ~n_24250 &  n_31218;
assign n_31220 = ~n_24244 &  n_31219;
assign n_31221 = ~n_24238 &  n_31220;
assign n_31222 = ~n_24232 &  n_31221;
assign n_31223 = ~n_24226 &  n_31222;
assign n_31224 = ~n_24219 &  n_31223;
assign n_31225 = ~n_24213 &  n_31224;
assign n_31226 = ~n_24207 &  n_31225;
assign n_31227 = ~n_24201 &  n_31226;
assign n_31228 = ~n_24195 &  n_31227;
assign n_31229 = ~n_24189 &  n_31228;
assign n_31230 = ~n_24183 &  n_31229;
assign n_31231 = ~n_24177 &  n_31230;
assign n_31232 = ~n_24171 &  n_31231;
assign n_31233 = ~n_24165 &  n_31232;
assign n_31234 = ~n_24159 &  n_31233;
assign n_31235 = ~n_24153 &  n_31234;
assign n_31236 = ~n_24147 &  n_31235;
assign n_31237 = ~n_24141 &  n_31236;
assign n_31238 = ~n_24135 &  n_31237;
assign n_31239 = ~n_24129 &  n_31238;
assign n_31240 = ~n_24123 &  n_31239;
assign n_31241 = ~n_24117 &  n_31240;
assign n_31242 = ~n_24111 &  n_31241;
assign n_31243 = ~n_24105 &  n_31242;
assign n_31244 = ~n_24099 &  n_31243;
assign n_31245 = ~n_24093 &  n_31244;
assign n_31246 = ~n_24087 &  n_31245;
assign n_31247 = ~n_24081 &  n_31246;
assign n_31248 = ~n_24075 &  n_31247;
assign n_31249 = ~n_24069 &  n_31248;
assign n_31250 = ~n_24063 &  n_31249;
assign n_31251 = ~n_24057 &  n_31250;
assign n_31252 = ~n_24051 &  n_31251;
assign n_31253 = ~n_24045 &  n_31252;
assign n_31254 = ~n_24039 &  n_31253;
assign n_31255 = ~n_24033 &  n_31254;
assign n_31256 = ~n_24026 &  n_31255;
assign n_31257 = ~n_24022 &  n_31256;
assign n_31258 = ~n_24018 &  n_31257;
assign n_31259 = ~n_24014 &  n_31258;
assign n_31260 = ~n_24010 &  n_31259;
assign n_31261 = ~n_24006 &  n_31260;
assign n_31262 = ~n_24002 &  n_31261;
assign n_31263 = ~n_23998 &  n_31262;
assign n_31264 = ~n_23994 &  n_31263;
assign n_31265 = ~n_23990 &  n_31264;
assign n_31266 = ~n_23986 &  n_31265;
assign n_31267 = ~n_23982 &  n_31266;
assign n_31268 = ~n_23978 &  n_31267;
assign n_31269 = ~n_23974 &  n_31268;
assign n_31270 = ~n_23970 &  n_31269;
assign n_31271 = ~n_23966 &  n_31270;
assign n_31272 = ~n_23962 &  n_31271;
assign n_31273 = ~n_23958 &  n_31272;
assign n_31274 = ~n_23954 &  n_31273;
assign n_31275 = ~n_23950 &  n_31274;
assign n_31276 = ~n_23946 &  n_31275;
assign n_31277 = ~n_23942 &  n_31276;
assign n_31278 = ~n_23938 &  n_31277;
assign n_31279 = ~n_23934 &  n_31278;
assign n_31280 = ~n_23930 &  n_31279;
assign n_31281 = ~n_23926 &  n_31280;
assign n_31282 = ~n_23922 &  n_31281;
assign n_31283 = ~n_23918 &  n_31282;
assign n_31284 = ~n_23914 &  n_31283;
assign n_31285 = ~n_23910 &  n_31284;
assign n_31286 = ~n_23906 &  n_31285;
assign n_31287 = ~n_23902 &  n_31286;
assign n_31288 = ~n_23890 &  n_31287;
assign n_31289 = ~n_23884 &  n_31288;
assign n_31290 = ~n_23878 &  n_31289;
assign n_31291 = ~n_23872 &  n_31290;
assign n_31292 = ~n_23866 &  n_31291;
assign n_31293 = ~n_23860 &  n_31292;
assign n_31294 = ~n_23854 &  n_31293;
assign n_31295 = ~n_23848 &  n_31294;
assign n_31296 = ~n_23842 &  n_31295;
assign n_31297 = ~n_23836 &  n_31296;
assign n_31298 = ~n_23830 &  n_31297;
assign n_31299 = ~n_23824 &  n_31298;
assign n_31300 = ~n_23818 &  n_31299;
assign n_31301 = ~n_23812 &  n_31300;
assign n_31302 = ~n_23806 &  n_31301;
assign n_31303 = ~n_23800 &  n_31302;
assign n_31304 = ~n_23794 &  n_31303;
assign n_31305 = ~n_23788 &  n_31304;
assign n_31306 = ~n_23782 &  n_31305;
assign n_31307 = ~n_23776 &  n_31306;
assign n_31308 = ~n_23770 &  n_31307;
assign n_31309 = ~n_23764 &  n_31308;
assign n_31310 = ~n_23758 &  n_31309;
assign n_31311 = ~n_23752 &  n_31310;
assign n_31312 = ~n_23746 &  n_31311;
assign n_31313 = ~n_23740 &  n_31312;
assign n_31314 = ~n_23734 &  n_31313;
assign n_31315 = ~n_23728 &  n_31314;
assign n_31316 = ~n_23722 &  n_31315;
assign n_31317 = ~n_23716 &  n_31316;
assign n_31318 = ~n_23710 &  n_31317;
assign n_31319 = ~n_23704 &  n_31318;
assign n_31320 = ~n_23696 &  n_31319;
assign n_31321 = ~n_23690 &  n_31320;
assign n_31322 = ~n_23684 &  n_31321;
assign n_31323 = ~n_23678 &  n_31322;
assign n_31324 = ~n_23672 &  n_31323;
assign n_31325 = ~n_23666 &  n_31324;
assign n_31326 = ~n_23660 &  n_31325;
assign n_31327 = ~n_23654 &  n_31326;
assign n_31328 = ~n_23648 &  n_31327;
assign n_31329 = ~n_23642 &  n_31328;
assign n_31330 = ~n_23636 &  n_31329;
assign n_31331 = ~n_23630 &  n_31330;
assign n_31332 = ~n_23624 &  n_31331;
assign n_31333 = ~n_23618 &  n_31332;
assign n_31334 = ~n_23612 &  n_31333;
assign n_31335 = ~n_23606 &  n_31334;
assign n_31336 = ~n_23600 &  n_31335;
assign n_31337 = ~n_23594 &  n_31336;
assign n_31338 = ~n_23588 &  n_31337;
assign n_31339 = ~n_23582 &  n_31338;
assign n_31340 = ~n_23576 &  n_31339;
assign n_31341 = ~n_23570 &  n_31340;
assign n_31342 = ~n_23564 &  n_31341;
assign n_31343 = ~n_23558 &  n_31342;
assign n_31344 = ~n_23552 &  n_31343;
assign n_31345 = ~n_23546 &  n_31344;
assign n_31346 = ~n_23540 &  n_31345;
assign n_31347 = ~n_23534 &  n_31346;
assign n_31348 = ~n_23528 &  n_31347;
assign n_31349 = ~n_23522 &  n_31348;
assign n_31350 = ~n_23516 &  n_31349;
assign n_31351 = ~n_23510 &  n_31350;
assign n_31352 = ~n_23502 &  n_31351;
assign n_31353 = ~n_23496 &  n_31352;
assign n_31354 = ~n_23490 &  n_31353;
assign n_31355 = ~n_23484 &  n_31354;
assign n_31356 = ~n_23478 &  n_31355;
assign n_31357 = ~n_23472 &  n_31356;
assign n_31358 = ~n_23466 &  n_31357;
assign n_31359 = ~n_23460 &  n_31358;
assign n_31360 = ~n_23454 &  n_31359;
assign n_31361 = ~n_23448 &  n_31360;
assign n_31362 = ~n_23442 &  n_31361;
assign n_31363 = ~n_23436 &  n_31362;
assign n_31364 = ~n_23430 &  n_31363;
assign n_31365 = ~n_23424 &  n_31364;
assign n_31366 = ~n_23418 &  n_31365;
assign n_31367 = ~n_23412 &  n_31366;
assign n_31368 = ~n_23406 &  n_31367;
assign n_31369 = ~n_23400 &  n_31368;
assign n_31370 = ~n_23394 &  n_31369;
assign n_31371 = ~n_23388 &  n_31370;
assign n_31372 = ~n_23382 &  n_31371;
assign n_31373 = ~n_23376 &  n_31372;
assign n_31374 = ~n_23370 &  n_31373;
assign n_31375 = ~n_23364 &  n_31374;
assign n_31376 = ~n_23358 &  n_31375;
assign n_31377 = ~n_23352 &  n_31376;
assign n_31378 = ~n_23346 &  n_31377;
assign n_31379 = ~n_23340 &  n_31378;
assign n_31380 = ~n_23334 &  n_31379;
assign n_31381 = ~n_23328 &  n_31380;
assign n_31382 = ~n_23322 &  n_31381;
assign n_31383 = ~n_23316 &  n_31382;
assign n_31384 = ~n_23309 &  n_31383;
assign n_31385 = ~n_23303 &  n_31384;
assign n_31386 = ~n_23297 &  n_31385;
assign n_31387 = ~n_23291 &  n_31386;
assign n_31388 = ~n_23285 &  n_31387;
assign n_31389 = ~n_23279 &  n_31388;
assign n_31390 = ~n_23273 &  n_31389;
assign n_31391 = ~n_23267 &  n_31390;
assign n_31392 = ~n_23261 &  n_31391;
assign n_31393 = ~n_23255 &  n_31392;
assign n_31394 = ~n_23249 &  n_31393;
assign n_31395 = ~n_23243 &  n_31394;
assign n_31396 = ~n_23237 &  n_31395;
assign n_31397 = ~n_23231 &  n_31396;
assign n_31398 = ~n_23225 &  n_31397;
assign n_31399 = ~n_23219 &  n_31398;
assign n_31400 = ~n_23213 &  n_31399;
assign n_31401 = ~n_23207 &  n_31400;
assign n_31402 = ~n_23201 &  n_31401;
assign n_31403 = ~n_23195 &  n_31402;
assign n_31404 = ~n_23189 &  n_31403;
assign n_31405 = ~n_23183 &  n_31404;
assign n_31406 = ~n_23177 &  n_31405;
assign n_31407 = ~n_23171 &  n_31406;
assign n_31408 = ~n_23165 &  n_31407;
assign n_31409 = ~n_23159 &  n_31408;
assign n_31410 = ~n_23153 &  n_31409;
assign n_31411 = ~n_23147 &  n_31410;
assign n_31412 = ~n_23141 &  n_31411;
assign n_31413 = ~n_23135 &  n_31412;
assign n_31414 = ~n_23129 &  n_31413;
assign n_31415 = ~n_23123 &  n_31414;
assign n_31416 = ~n_23116 &  n_31415;
assign n_31417 = ~n_23110 &  n_31416;
assign n_31418 = ~n_23104 &  n_31417;
assign n_31419 = ~n_23098 &  n_31418;
assign n_31420 = ~n_23092 &  n_31419;
assign n_31421 = ~n_23086 &  n_31420;
assign n_31422 = ~n_23080 &  n_31421;
assign n_31423 = ~n_23074 &  n_31422;
assign n_31424 = ~n_23068 &  n_31423;
assign n_31425 = ~n_23062 &  n_31424;
assign n_31426 = ~n_23056 &  n_31425;
assign n_31427 = ~n_23050 &  n_31426;
assign n_31428 = ~n_23044 &  n_31427;
assign n_31429 = ~n_23038 &  n_31428;
assign n_31430 = ~n_23032 &  n_31429;
assign n_31431 = ~n_23026 &  n_31430;
assign n_31432 = ~n_23020 &  n_31431;
assign n_31433 = ~n_23014 &  n_31432;
assign n_31434 = ~n_23008 &  n_31433;
assign n_31435 = ~n_23002 &  n_31434;
assign n_31436 = ~n_22996 &  n_31435;
assign n_31437 = ~n_22990 &  n_31436;
assign n_31438 = ~n_22984 &  n_31437;
assign n_31439 = ~n_22978 &  n_31438;
assign n_31440 = ~n_22972 &  n_31439;
assign n_31441 = ~n_22966 &  n_31440;
assign n_31442 = ~n_22960 &  n_31441;
assign n_31443 = ~n_22954 &  n_31442;
assign n_31444 = ~n_22948 &  n_31443;
assign n_31445 = ~n_22942 &  n_31444;
assign n_31446 = ~n_22936 &  n_31445;
assign n_31447 = ~n_22930 &  n_31446;
assign n_31448 = ~n_22923 &  n_31447;
assign n_31449 = ~n_22917 &  n_31448;
assign n_31450 = ~n_22911 &  n_31449;
assign n_31451 = ~n_22905 &  n_31450;
assign n_31452 = ~n_22899 &  n_31451;
assign n_31453 = ~n_22893 &  n_31452;
assign n_31454 = ~n_22887 &  n_31453;
assign n_31455 = ~n_22881 &  n_31454;
assign n_31456 = ~n_22875 &  n_31455;
assign n_31457 = ~n_22869 &  n_31456;
assign n_31458 = ~n_22863 &  n_31457;
assign n_31459 = ~n_22857 &  n_31458;
assign n_31460 = ~n_22851 &  n_31459;
assign n_31461 = ~n_22845 &  n_31460;
assign n_31462 = ~n_22839 &  n_31461;
assign n_31463 = ~n_22833 &  n_31462;
assign n_31464 = ~n_22827 &  n_31463;
assign n_31465 = ~n_22821 &  n_31464;
assign n_31466 = ~n_22815 &  n_31465;
assign n_31467 = ~n_22809 &  n_31466;
assign n_31468 = ~n_22803 &  n_31467;
assign n_31469 = ~n_22797 &  n_31468;
assign n_31470 = ~n_22791 &  n_31469;
assign n_31471 = ~n_22785 &  n_31470;
assign n_31472 = ~n_22779 &  n_31471;
assign n_31473 = ~n_22773 &  n_31472;
assign n_31474 = ~n_22767 &  n_31473;
assign n_31475 = ~n_22761 &  n_31474;
assign n_31476 = ~n_22755 &  n_31475;
assign n_31477 = ~n_22749 &  n_31476;
assign n_31478 = ~n_22743 &  n_31477;
assign n_31479 = ~n_22737 &  n_31478;
assign n_31480 = ~n_22730 &  n_31479;
assign n_31481 = ~n_22724 &  n_31480;
assign n_31482 = ~n_22718 &  n_31481;
assign n_31483 = ~n_22712 &  n_31482;
assign n_31484 = ~n_22706 &  n_31483;
assign n_31485 = ~n_22700 &  n_31484;
assign n_31486 = ~n_22694 &  n_31485;
assign n_31487 = ~n_22688 &  n_31486;
assign n_31488 = ~n_22682 &  n_31487;
assign n_31489 = ~n_22676 &  n_31488;
assign n_31490 = ~n_22670 &  n_31489;
assign n_31491 = ~n_22664 &  n_31490;
assign n_31492 = ~n_22658 &  n_31491;
assign n_31493 = ~n_22652 &  n_31492;
assign n_31494 = ~n_22646 &  n_31493;
assign n_31495 = ~n_22640 &  n_31494;
assign n_31496 = ~n_22634 &  n_31495;
assign n_31497 = ~n_22628 &  n_31496;
assign n_31498 = ~n_22622 &  n_31497;
assign n_31499 = ~n_22616 &  n_31498;
assign n_31500 = ~n_22610 &  n_31499;
assign n_31501 = ~n_22604 &  n_31500;
assign n_31502 = ~n_22598 &  n_31501;
assign n_31503 = ~n_22592 &  n_31502;
assign n_31504 = ~n_22586 &  n_31503;
assign n_31505 = ~n_22580 &  n_31504;
assign n_31506 = ~n_22574 &  n_31505;
assign n_31507 = ~n_22568 &  n_31506;
assign n_31508 = ~n_22562 &  n_31507;
assign n_31509 = ~n_22556 &  n_31508;
assign n_31510 = ~n_22550 &  n_31509;
assign n_31511 = ~n_22544 &  n_31510;
assign n_31512 = ~n_22537 &  n_31511;
assign n_31513 = ~n_22531 &  n_31512;
assign n_31514 = ~n_22525 &  n_31513;
assign n_31515 = ~n_22519 &  n_31514;
assign n_31516 = ~n_22513 &  n_31515;
assign n_31517 = ~n_22507 &  n_31516;
assign n_31518 = ~n_22501 &  n_31517;
assign n_31519 = ~n_22495 &  n_31518;
assign n_31520 = ~n_22489 &  n_31519;
assign n_31521 = ~n_22483 &  n_31520;
assign n_31522 = ~n_22477 &  n_31521;
assign n_31523 = ~n_22471 &  n_31522;
assign n_31524 = ~n_22465 &  n_31523;
assign n_31525 = ~n_22459 &  n_31524;
assign n_31526 = ~n_22453 &  n_31525;
assign n_31527 = ~n_22447 &  n_31526;
assign n_31528 = ~n_22441 &  n_31527;
assign n_31529 = ~n_22435 &  n_31528;
assign n_31530 = ~n_22429 &  n_31529;
assign n_31531 = ~n_22423 &  n_31530;
assign n_31532 = ~n_22417 &  n_31531;
assign n_31533 = ~n_22411 &  n_31532;
assign n_31534 = ~n_22405 &  n_31533;
assign n_31535 = ~n_22399 &  n_31534;
assign n_31536 = ~n_22393 &  n_31535;
assign n_31537 = ~n_22387 &  n_31536;
assign n_31538 = ~n_22381 &  n_31537;
assign n_31539 = ~n_22375 &  n_31538;
assign n_31540 = ~n_22369 &  n_31539;
assign n_31541 = ~n_22363 &  n_31540;
assign n_31542 = ~n_22357 &  n_31541;
assign n_31543 = ~n_22351 &  n_31542;
assign n_31544 = ~n_22344 &  n_31543;
assign n_31545 = ~n_22338 &  n_31544;
assign n_31546 = ~n_22332 &  n_31545;
assign n_31547 = ~n_22326 &  n_31546;
assign n_31548 = ~n_22320 &  n_31547;
assign n_31549 = ~n_22314 &  n_31548;
assign n_31550 = ~n_22308 &  n_31549;
assign n_31551 = ~n_22302 &  n_31550;
assign n_31552 = ~n_22296 &  n_31551;
assign n_31553 = ~n_22290 &  n_31552;
assign n_31554 = ~n_22284 &  n_31553;
assign n_31555 = ~n_22278 &  n_31554;
assign n_31556 = ~n_22272 &  n_31555;
assign n_31557 = ~n_22264 &  n_31556;
assign n_31558 = ~n_22258 &  n_31557;
assign n_31559 = ~n_22252 &  n_31558;
assign n_31560 = ~n_22246 &  n_31559;
assign n_31561 = ~n_22240 &  n_31560;
assign n_31562 = ~n_22234 &  n_31561;
assign n_31563 = ~n_22228 &  n_31562;
assign n_31564 = ~n_22222 &  n_31563;
assign n_31565 = ~n_22216 &  n_31564;
assign n_31566 = ~n_22210 &  n_31565;
assign n_31567 = ~n_22204 &  n_31566;
assign n_31568 = ~n_22198 &  n_31567;
assign n_31569 = ~n_22192 &  n_31568;
assign n_31570 = ~n_22186 &  n_31569;
assign n_31571 = ~n_22180 &  n_31570;
assign n_31572 = ~n_22174 &  n_31571;
assign n_31573 = ~n_22168 &  n_31572;
assign n_31574 = ~n_22162 &  n_31573;
assign n_31575 = ~n_22156 &  n_31574;
assign n_31576 = ~n_22150 &  n_31575;
assign n_31577 = ~n_22144 &  n_31576;
assign n_31578 = ~n_22138 &  n_31577;
assign n_31579 = ~n_22132 &  n_31578;
assign n_31580 = ~n_22126 &  n_31579;
assign n_31581 = ~n_22120 &  n_31580;
assign n_31582 = ~n_22114 &  n_31581;
assign n_31583 = ~n_22108 &  n_31582;
assign n_31584 = ~n_22102 &  n_31583;
assign n_31585 = ~n_22096 &  n_31584;
assign n_31586 = ~n_22090 &  n_31585;
assign n_31587 = ~n_22084 &  n_31586;
assign n_31588 = ~n_22078 &  n_31587;
assign n_31589 = ~n_22071 &  n_31588;
assign n_31590 = ~n_22065 &  n_31589;
assign n_31591 = ~n_22059 &  n_31590;
assign n_31592 = ~n_22053 &  n_31591;
assign n_31593 = ~n_22047 &  n_31592;
assign n_31594 = ~n_22041 &  n_31593;
assign n_31595 = ~n_22035 &  n_31594;
assign n_31596 = ~n_22029 &  n_31595;
assign n_31597 = ~n_22023 &  n_31596;
assign n_31598 = ~n_22017 &  n_31597;
assign n_31599 = ~n_22011 &  n_31598;
assign n_31600 = ~n_22005 &  n_31599;
assign n_31601 = ~n_21999 &  n_31600;
assign n_31602 = ~n_21993 &  n_31601;
assign n_31603 = ~n_21987 &  n_31602;
assign n_31604 = ~n_21981 &  n_31603;
assign n_31605 = ~n_21975 &  n_31604;
assign n_31606 = ~n_21969 &  n_31605;
assign n_31607 = ~n_21963 &  n_31606;
assign n_31608 = ~n_21957 &  n_31607;
assign n_31609 = ~n_21951 &  n_31608;
assign n_31610 = ~n_21945 &  n_31609;
assign n_31611 = ~n_21939 &  n_31610;
assign n_31612 = ~n_21933 &  n_31611;
assign n_31613 = ~n_21927 &  n_31612;
assign n_31614 = ~n_21921 &  n_31613;
assign n_31615 = ~n_21915 &  n_31614;
assign n_31616 = ~n_21909 &  n_31615;
assign n_31617 = ~n_21903 &  n_31616;
assign n_31618 = ~n_21897 &  n_31617;
assign n_31619 = ~n_21891 &  n_31618;
assign n_31620 = ~n_21885 &  n_31619;
assign n_31621 = ~n_21878 &  n_31620;
assign n_31622 = ~n_21872 &  n_31621;
assign n_31623 = ~n_21866 &  n_31622;
assign n_31624 = ~n_21860 &  n_31623;
assign n_31625 = ~n_21854 &  n_31624;
assign n_31626 = ~n_21848 &  n_31625;
assign n_31627 = ~n_21842 &  n_31626;
assign n_31628 = ~n_21836 &  n_31627;
assign n_31629 = ~n_21830 &  n_31628;
assign n_31630 = ~n_21824 &  n_31629;
assign n_31631 = ~n_21818 &  n_31630;
assign n_31632 = ~n_21812 &  n_31631;
assign n_31633 = ~n_21806 &  n_31632;
assign n_31634 = ~n_21800 &  n_31633;
assign n_31635 = ~n_21794 &  n_31634;
assign n_31636 = ~n_21788 &  n_31635;
assign n_31637 = ~n_21782 &  n_31636;
assign n_31638 = ~n_21776 &  n_31637;
assign n_31639 = ~n_21770 &  n_31638;
assign n_31640 = ~n_21764 &  n_31639;
assign n_31641 = ~n_21758 &  n_31640;
assign n_31642 = ~n_21752 &  n_31641;
assign n_31643 = ~n_21746 &  n_31642;
assign n_31644 = ~n_21740 &  n_31643;
assign n_31645 = ~n_21734 &  n_31644;
assign n_31646 = ~n_21728 &  n_31645;
assign n_31647 = ~n_21722 &  n_31646;
assign n_31648 = ~n_21716 &  n_31647;
assign n_31649 = ~n_21710 &  n_31648;
assign n_31650 = ~n_21704 &  n_31649;
assign n_31651 = ~n_21698 &  n_31650;
assign n_31652 = ~n_21692 &  n_31651;
assign n_31653 = ~n_21685 &  n_31652;
assign n_31654 = ~n_21679 &  n_31653;
assign n_31655 = ~n_21673 &  n_31654;
assign n_31656 = ~n_21667 &  n_31655;
assign n_31657 = ~n_21661 &  n_31656;
assign n_31658 = ~n_21655 &  n_31657;
assign n_31659 = ~n_21649 &  n_31658;
assign n_31660 = ~n_21643 &  n_31659;
assign n_31661 = ~n_21637 &  n_31660;
assign n_31662 = ~n_21631 &  n_31661;
assign n_31663 = ~n_21625 &  n_31662;
assign n_31664 = ~n_21619 &  n_31663;
assign n_31665 = ~n_21613 &  n_31664;
assign n_31666 = ~n_21607 &  n_31665;
assign n_31667 = ~n_21601 &  n_31666;
assign n_31668 = ~n_21595 &  n_31667;
assign n_31669 = ~n_21589 &  n_31668;
assign n_31670 = ~n_21583 &  n_31669;
assign n_31671 = ~n_21577 &  n_31670;
assign n_31672 = ~n_21571 &  n_31671;
assign n_31673 = ~n_21565 &  n_31672;
assign n_31674 = ~n_21559 &  n_31673;
assign n_31675 = ~n_21553 &  n_31674;
assign n_31676 = ~n_21547 &  n_31675;
assign n_31677 = ~n_21541 &  n_31676;
assign n_31678 = ~n_21535 &  n_31677;
assign n_31679 = ~n_21529 &  n_31678;
assign n_31680 = ~n_21523 &  n_31679;
assign n_31681 = ~n_21517 &  n_31680;
assign n_31682 = ~n_21511 &  n_31681;
assign n_31683 = ~n_21505 &  n_31682;
assign n_31684 = ~n_21499 &  n_31683;
assign n_31685 = ~n_21492 &  n_31684;
assign n_31686 = ~n_21486 &  n_31685;
assign n_31687 = ~n_21480 &  n_31686;
assign n_31688 = ~n_21474 &  n_31687;
assign n_31689 = ~n_21468 &  n_31688;
assign n_31690 = ~n_21462 &  n_31689;
assign n_31691 = ~n_21456 &  n_31690;
assign n_31692 = ~n_21450 &  n_31691;
assign n_31693 = ~n_21444 &  n_31692;
assign n_31694 = ~n_21438 &  n_31693;
assign n_31695 = ~n_21432 &  n_31694;
assign n_31696 = ~n_21426 &  n_31695;
assign n_31697 = ~n_21420 &  n_31696;
assign n_31698 = ~n_21414 &  n_31697;
assign n_31699 = ~n_21408 &  n_31698;
assign n_31700 = ~n_21402 &  n_31699;
assign n_31701 = ~n_21396 &  n_31700;
assign n_31702 = ~n_21390 &  n_31701;
assign n_31703 = ~n_21384 &  n_31702;
assign n_31704 = ~n_21378 &  n_31703;
assign n_31705 = ~n_21372 &  n_31704;
assign n_31706 = ~n_21366 &  n_31705;
assign n_31707 = ~n_21360 &  n_31706;
assign n_31708 = ~n_21354 &  n_31707;
assign n_31709 = ~n_21348 &  n_31708;
assign n_31710 = ~n_21342 &  n_31709;
assign n_31711 = ~n_21336 &  n_31710;
assign n_31712 = ~n_21330 &  n_31711;
assign n_31713 = ~n_21324 &  n_31712;
assign n_31714 = ~n_21318 &  n_31713;
assign n_31715 = ~n_21312 &  n_31714;
assign n_31716 = ~n_21306 &  n_31715;
assign n_31717 = ~n_21299 &  n_31716;
assign n_31718 = ~n_21293 &  n_31717;
assign n_31719 = ~n_21287 &  n_31718;
assign n_31720 = ~n_21281 &  n_31719;
assign n_31721 = ~n_21275 &  n_31720;
assign n_31722 = ~n_21269 &  n_31721;
assign n_31723 = ~n_21263 &  n_31722;
assign n_31724 = ~n_21257 &  n_31723;
assign n_31725 = ~n_21251 &  n_31724;
assign n_31726 = ~n_21245 &  n_31725;
assign n_31727 = ~n_21239 &  n_31726;
assign n_31728 = ~n_21233 &  n_31727;
assign n_31729 = ~n_21227 &  n_31728;
assign n_31730 = ~n_21221 &  n_31729;
assign n_31731 = ~n_21215 &  n_31730;
assign n_31732 = ~n_21209 &  n_31731;
assign n_31733 = ~n_21203 &  n_31732;
assign n_31734 = ~n_21197 &  n_31733;
assign n_31735 = ~n_21191 &  n_31734;
assign n_31736 = ~n_21185 &  n_31735;
assign n_31737 = ~n_21179 &  n_31736;
assign n_31738 = ~n_21173 &  n_31737;
assign n_31739 = ~n_21167 &  n_31738;
assign n_31740 = ~n_21161 &  n_31739;
assign n_31741 = ~n_21155 &  n_31740;
assign n_31742 = ~n_21149 &  n_31741;
assign n_31743 = ~n_21143 &  n_31742;
assign n_31744 = ~n_21137 &  n_31743;
assign n_31745 = ~n_21131 &  n_31744;
assign n_31746 = ~n_21125 &  n_31745;
assign n_31747 = ~n_21119 &  n_31746;
assign n_31748 = ~n_21113 &  n_31747;
assign n_31749 = ~n_21106 &  n_31748;
assign n_31750 = ~n_21100 &  n_31749;
assign n_31751 = ~n_21094 &  n_31750;
assign n_31752 = ~n_21088 &  n_31751;
assign n_31753 = ~n_21082 &  n_31752;
assign n_31754 = ~n_21076 &  n_31753;
assign n_31755 = ~n_21070 &  n_31754;
assign n_31756 = ~n_21064 &  n_31755;
assign n_31757 = ~n_21058 &  n_31756;
assign n_31758 = ~n_21052 &  n_31757;
assign n_31759 = ~n_21046 &  n_31758;
assign n_31760 = ~n_21040 &  n_31759;
assign n_31761 = ~n_21034 &  n_31760;
assign n_31762 = ~n_21028 &  n_31761;
assign n_31763 = ~n_21022 &  n_31762;
assign n_31764 = ~n_21016 &  n_31763;
assign n_31765 = ~n_21010 &  n_31764;
assign n_31766 = ~n_21004 &  n_31765;
assign n_31767 = ~n_20998 &  n_31766;
assign n_31768 = ~n_20992 &  n_31767;
assign n_31769 = ~n_20986 &  n_31768;
assign n_31770 = ~n_20980 &  n_31769;
assign n_31771 = ~n_20974 &  n_31770;
assign n_31772 = ~n_20968 &  n_31771;
assign n_31773 = ~n_20962 &  n_31772;
assign n_31774 = ~n_20956 &  n_31773;
assign n_31775 = ~n_20950 &  n_31774;
assign n_31776 = ~n_20944 &  n_31775;
assign n_31777 = ~n_20938 &  n_31776;
assign n_31778 = ~n_20932 &  n_31777;
assign n_31779 = ~n_20926 &  n_31778;
assign n_31780 = ~n_20920 &  n_31779;
assign n_31781 = ~n_20913 &  n_31780;
assign n_31782 = ~n_20907 &  n_31781;
assign n_31783 = ~n_20901 &  n_31782;
assign n_31784 = ~n_20895 &  n_31783;
assign n_31785 = ~n_20889 &  n_31784;
assign n_31786 = ~n_20883 &  n_31785;
assign n_31787 = ~n_20877 &  n_31786;
assign n_31788 = ~n_20871 &  n_31787;
assign n_31789 = ~n_20865 &  n_31788;
assign n_31790 = ~n_20859 &  n_31789;
assign n_31791 = ~n_20853 &  n_31790;
assign n_31792 = ~n_20847 &  n_31791;
assign n_31793 = ~n_20841 &  n_31792;
assign n_31794 = ~n_20835 &  n_31793;
assign n_31795 = ~n_20829 &  n_31794;
assign n_31796 = ~n_20823 &  n_31795;
assign n_31797 = ~n_20817 &  n_31796;
assign n_31798 = ~n_20811 &  n_31797;
assign n_31799 = ~n_20805 &  n_31798;
assign n_31800 = ~n_20799 &  n_31799;
assign n_31801 = ~n_20793 &  n_31800;
assign n_31802 = ~n_20787 &  n_31801;
assign n_31803 = ~n_20781 &  n_31802;
assign n_31804 = ~n_20775 &  n_31803;
assign n_31805 = ~n_20769 &  n_31804;
assign n_31806 = ~n_20763 &  n_31805;
assign n_31807 = ~n_20757 &  n_31806;
assign n_31808 = ~n_20751 &  n_31807;
assign n_31809 = ~n_20745 &  n_31808;
assign n_31810 = ~n_20739 &  n_31809;
assign n_31811 = ~n_20733 &  n_31810;
assign n_31812 = ~n_20727 &  n_31811;
assign n_31813 = ~n_20717 &  n_31812;
assign n_31814 = ~n_20711 &  n_31813;
assign n_31815 = ~n_20705 &  n_31814;
assign n_31816 = ~n_20699 &  n_31815;
assign n_31817 = ~n_20693 &  n_31816;
assign n_31818 = ~n_20687 &  n_31817;
assign n_31819 = ~n_20681 &  n_31818;
assign n_31820 = ~n_20675 &  n_31819;
assign n_31821 = ~n_20669 &  n_31820;
assign n_31822 = ~n_20663 &  n_31821;
assign n_31823 = ~n_20657 &  n_31822;
assign n_31824 = ~n_20651 &  n_31823;
assign n_31825 = ~n_20645 &  n_31824;
assign n_31826 = ~n_20639 &  n_31825;
assign n_31827 = ~n_20633 &  n_31826;
assign n_31828 = ~n_20627 &  n_31827;
assign n_31829 = ~n_20621 &  n_31828;
assign n_31830 = ~n_20615 &  n_31829;
assign n_31831 = ~n_20609 &  n_31830;
assign n_31832 = ~n_20603 &  n_31831;
assign n_31833 = ~n_20597 &  n_31832;
assign n_31834 = ~n_20591 &  n_31833;
assign n_31835 = ~n_20585 &  n_31834;
assign n_31836 = ~n_20579 &  n_31835;
assign n_31837 = ~n_20573 &  n_31836;
assign n_31838 = ~n_20567 &  n_31837;
assign n_31839 = ~n_20561 &  n_31838;
assign n_31840 = ~n_20555 &  n_31839;
assign n_31841 = ~n_20549 &  n_31840;
assign n_31842 = ~n_20543 &  n_31841;
assign n_31843 = ~n_20537 &  n_31842;
assign n_31844 = ~n_20531 &  n_31843;
assign n_31845 = ~n_20524 &  n_31844;
assign n_31846 = ~n_20518 &  n_31845;
assign n_31847 = ~n_20512 &  n_31846;
assign n_31848 = ~n_20506 &  n_31847;
assign n_31849 = ~n_20500 &  n_31848;
assign n_31850 = ~n_20494 &  n_31849;
assign n_31851 = ~n_20488 &  n_31850;
assign n_31852 = ~n_20482 &  n_31851;
assign n_31853 = ~n_20476 &  n_31852;
assign n_31854 = ~n_20470 &  n_31853;
assign n_31855 = ~n_20464 &  n_31854;
assign n_31856 = ~n_20458 &  n_31855;
assign n_31857 = ~n_20452 &  n_31856;
assign n_31858 = ~n_20446 &  n_31857;
assign n_31859 = ~n_20440 &  n_31858;
assign n_31860 = ~n_20434 &  n_31859;
assign n_31861 = ~n_20428 &  n_31860;
assign n_31862 = ~n_20422 &  n_31861;
assign n_31863 = ~n_20416 &  n_31862;
assign n_31864 = ~n_20410 &  n_31863;
assign n_31865 = ~n_20404 &  n_31864;
assign n_31866 = ~n_20398 &  n_31865;
assign n_31867 = ~n_20392 &  n_31866;
assign n_31868 = ~n_20386 &  n_31867;
assign n_31869 = ~n_20380 &  n_31868;
assign n_31870 = ~n_20374 &  n_31869;
assign n_31871 = ~n_20368 &  n_31870;
assign n_31872 = ~n_20362 &  n_31871;
assign n_31873 = ~n_20356 &  n_31872;
assign n_31874 = ~n_20350 &  n_31873;
assign n_31875 = ~n_20344 &  n_31874;
assign n_31876 = ~n_20338 &  n_31875;
assign n_31877 = ~n_20331 &  n_31876;
assign n_31878 = ~n_20325 &  n_31877;
assign n_31879 = ~n_20319 &  n_31878;
assign n_31880 = ~n_20313 &  n_31879;
assign n_31881 = ~n_20307 &  n_31880;
assign n_31882 = ~n_20301 &  n_31881;
assign n_31883 = ~n_20295 &  n_31882;
assign n_31884 = ~n_20289 &  n_31883;
assign n_31885 = ~n_20283 &  n_31884;
assign n_31886 = ~n_20277 &  n_31885;
assign n_31887 = ~n_20271 &  n_31886;
assign n_31888 = ~n_20265 &  n_31887;
assign n_31889 = ~n_20259 &  n_31888;
assign n_31890 = ~n_20253 &  n_31889;
assign n_31891 = ~n_20247 &  n_31890;
assign n_31892 = ~n_20241 &  n_31891;
assign n_31893 = ~n_20235 &  n_31892;
assign n_31894 = ~n_20229 &  n_31893;
assign n_31895 = ~n_20223 &  n_31894;
assign n_31896 = ~n_20217 &  n_31895;
assign n_31897 = ~n_20211 &  n_31896;
assign n_31898 = ~n_20205 &  n_31897;
assign n_31899 = ~n_20199 &  n_31898;
assign n_31900 = ~n_20193 &  n_31899;
assign n_31901 = ~n_20187 &  n_31900;
assign n_31902 = ~n_20181 &  n_31901;
assign n_31903 = ~n_20175 &  n_31902;
assign n_31904 = ~n_20169 &  n_31903;
assign n_31905 = ~n_20163 &  n_31904;
assign n_31906 = ~n_20157 &  n_31905;
assign n_31907 = ~n_20151 &  n_31906;
assign n_31908 = ~n_20145 &  n_31907;
assign n_31909 = ~n_20138 &  n_31908;
assign n_31910 = ~n_20132 &  n_31909;
assign n_31911 = ~n_20126 &  n_31910;
assign n_31912 = ~n_20120 &  n_31911;
assign n_31913 = ~n_20114 &  n_31912;
assign n_31914 = ~n_20108 &  n_31913;
assign n_31915 = ~n_20102 &  n_31914;
assign n_31916 = ~n_20096 &  n_31915;
assign n_31917 = ~n_20090 &  n_31916;
assign n_31918 = ~n_20084 &  n_31917;
assign n_31919 = ~n_20078 &  n_31918;
assign n_31920 = ~n_20072 &  n_31919;
assign n_31921 = ~n_20066 &  n_31920;
assign n_31922 = ~n_20060 &  n_31921;
assign n_31923 = ~n_20054 &  n_31922;
assign n_31924 = ~n_20048 &  n_31923;
assign n_31925 = ~n_20042 &  n_31924;
assign n_31926 = ~n_20036 &  n_31925;
assign n_31927 = ~n_20030 &  n_31926;
assign n_31928 = ~n_20024 &  n_31927;
assign n_31929 = ~n_20018 &  n_31928;
assign n_31930 = ~n_20012 &  n_31929;
assign n_31931 = ~n_20006 &  n_31930;
assign n_31932 = ~n_20000 &  n_31931;
assign n_31933 = ~n_19994 &  n_31932;
assign n_31934 = ~n_19988 &  n_31933;
assign n_31935 = ~n_19982 &  n_31934;
assign n_31936 = ~n_19976 &  n_31935;
assign n_31937 = ~n_19970 &  n_31936;
assign n_31938 = ~n_19964 &  n_31937;
assign n_31939 = ~n_19958 &  n_31938;
assign n_31940 = ~n_19952 &  n_31939;
assign n_31941 = ~n_19944 &  n_31940;
assign n_31942 = ~n_19898 &  n_31941;
assign n_31943 = ~n_19850 &  n_31942;
assign n_31944 = ~n_19802 &  n_31943;
assign n_31945 = ~n_19754 &  n_31944;
assign n_31946 = ~n_19706 &  n_31945;
assign n_31947 = ~n_19658 &  n_31946;
assign n_31948 = ~n_19610 &  n_31947;
assign n_31949 = ~n_19562 &  n_31948;
assign n_31950 = ~n_19514 &  n_31949;
assign n_31951 = ~n_19466 &  n_31950;
assign n_31952 = ~n_19418 &  n_31951;
assign n_31953 = ~n_19370 &  n_31952;
assign n_31954 = ~n_19322 &  n_31953;
assign n_31955 = ~n_19274 &  n_31954;
assign n_31956 = ~n_19226 &  n_31955;
assign n_31957 = ~n_19178 &  n_31956;
assign n_31958 = ~n_19130 &  n_31957;
assign n_31959 = ~n_19082 &  n_31958;
assign n_31960 = ~n_19034 &  n_31959;
assign n_31961 = ~n_18986 &  n_31960;
assign n_31962 = ~n_18938 &  n_31961;
assign n_31963 = ~n_18890 &  n_31962;
assign n_31964 = ~n_18842 &  n_31963;
assign n_31965 = ~n_18794 &  n_31964;
assign n_31966 = ~n_18746 &  n_31965;
assign n_31967 = ~n_18698 &  n_31966;
assign n_31968 = ~n_18650 &  n_31967;
assign n_31969 = ~n_18602 &  n_31968;
assign n_31970 = ~n_18555 &  n_31969;
assign n_31971 = ~n_18501 &  n_31970;
assign n_31972 = ~n_18459 &  n_31971;
assign n_31973 = ~n_18428 &  n_31972;
assign n_31974 = ~n_18383 &  n_31973;
assign n_31975 = ~n_18335 &  n_31974;
assign n_31976 = ~n_18287 &  n_31975;
assign n_31977 = ~n_18239 &  n_31976;
assign n_31978 = ~n_18191 &  n_31977;
assign n_31979 = ~n_18143 &  n_31978;
assign n_31980 = ~n_18095 &  n_31979;
assign n_31981 = ~n_18047 &  n_31980;
assign n_31982 = ~n_17999 &  n_31981;
assign n_31983 = ~n_17951 &  n_31982;
assign n_31984 = ~n_17903 &  n_31983;
assign n_31985 = ~n_17855 &  n_31984;
assign n_31986 = ~n_17807 &  n_31985;
assign n_31987 = ~n_17759 &  n_31986;
assign n_31988 = ~n_17711 &  n_31987;
assign n_31989 = ~n_17663 &  n_31988;
assign n_31990 = ~n_17615 &  n_31989;
assign n_31991 = ~n_17567 &  n_31990;
assign n_31992 = ~n_17519 &  n_31991;
assign n_31993 = ~n_17471 &  n_31992;
assign n_31994 = ~n_17423 &  n_31993;
assign n_31995 = ~n_17375 &  n_31994;
assign n_31996 = ~n_17327 &  n_31995;
assign n_31997 = ~n_17279 &  n_31996;
assign n_31998 = ~n_17231 &  n_31997;
assign n_31999 = ~n_17183 &  n_31998;
assign n_32000 = ~n_17135 &  n_31999;
assign n_32001 = ~n_17087 &  n_32000;
assign n_32002 = ~n_17039 &  n_32001;
assign n_32003 = ~n_16985 &  n_32002;
assign n_32004 = ~n_16943 &  n_32003;
assign n_32005 = ~n_16913 &  n_32004;
assign n_32006 = ~n_16907 &  n_32005;
assign n_32007 = ~n_16901 &  n_32006;
assign n_32008 = ~n_16895 &  n_32007;
assign n_32009 = ~n_16889 &  n_32008;
assign n_32010 = ~n_16883 &  n_32009;
assign n_32011 = ~n_16877 &  n_32010;
assign n_32012 = ~n_16871 &  n_32011;
assign n_32013 = ~n_16865 &  n_32012;
assign n_32014 = ~n_16859 &  n_32013;
assign n_32015 = ~n_16853 &  n_32014;
assign n_32016 = ~n_16847 &  n_32015;
assign n_32017 = ~n_16841 &  n_32016;
assign n_32018 = ~n_16835 &  n_32017;
assign n_32019 = ~n_16829 &  n_32018;
assign n_32020 = ~n_16823 &  n_32019;
assign n_32021 = ~n_16817 &  n_32020;
assign n_32022 = ~n_16811 &  n_32021;
assign n_32023 = ~n_16805 &  n_32022;
assign n_32024 = ~n_16799 &  n_32023;
assign n_32025 = ~n_16793 &  n_32024;
assign n_32026 = ~n_16787 &  n_32025;
assign n_32027 = ~n_16781 &  n_32026;
assign n_32028 = ~n_16775 &  n_32027;
assign n_32029 = ~n_16769 &  n_32028;
assign n_32030 = ~n_16763 &  n_32029;
assign n_32031 = ~n_16757 &  n_32030;
assign n_32032 = ~n_16751 &  n_32031;
assign n_32033 = ~n_16745 &  n_32032;
assign n_32034 = ~n_16739 &  n_32033;
assign n_32035 = ~n_16733 &  n_32034;
assign n_32036 = ~n_16727 &  n_32035;
assign n_32037 = ~n_16720 &  n_32036;
assign n_32038 = ~n_16714 &  n_32037;
assign n_32039 = ~n_16708 &  n_32038;
assign n_32040 = ~n_16702 &  n_32039;
assign n_32041 = ~n_16696 &  n_32040;
assign n_32042 = ~n_16690 &  n_32041;
assign n_32043 = ~n_16684 &  n_32042;
assign n_32044 = ~n_16678 &  n_32043;
assign n_32045 = ~n_16672 &  n_32044;
assign n_32046 = ~n_16666 &  n_32045;
assign n_32047 = ~n_16660 &  n_32046;
assign n_32048 = ~n_16654 &  n_32047;
assign n_32049 = ~n_16648 &  n_32048;
assign n_32050 = ~n_16642 &  n_32049;
assign n_32051 = ~n_16636 &  n_32050;
assign n_32052 = ~n_16630 &  n_32051;
assign n_32053 = ~n_16624 &  n_32052;
assign n_32054 = ~n_16618 &  n_32053;
assign n_32055 = ~n_16612 &  n_32054;
assign n_32056 = ~n_16606 &  n_32055;
assign n_32057 = ~n_16600 &  n_32056;
assign n_32058 = ~n_16594 &  n_32057;
assign n_32059 = ~n_16588 &  n_32058;
assign n_32060 = ~n_16582 &  n_32059;
assign n_32061 = ~n_16576 &  n_32060;
assign n_32062 = ~n_16570 &  n_32061;
assign n_32063 = ~n_16564 &  n_32062;
assign n_32064 = ~n_16558 &  n_32063;
assign n_32065 = ~n_16552 &  n_32064;
assign n_32066 = ~n_16546 &  n_32065;
assign n_32067 = ~n_16540 &  n_32066;
assign n_32068 = ~n_16534 &  n_32067;
assign n_32069 = ~n_16527 &  n_32068;
assign n_32070 = ~n_16521 &  n_32069;
assign n_32071 = ~n_16515 &  n_32070;
assign n_32072 = ~n_16509 &  n_32071;
assign n_32073 = ~n_16503 &  n_32072;
assign n_32074 = ~n_16497 &  n_32073;
assign n_32075 = ~n_16491 &  n_32074;
assign n_32076 = ~n_16485 &  n_32075;
assign n_32077 = ~n_16479 &  n_32076;
assign n_32078 = ~n_16473 &  n_32077;
assign n_32079 = ~n_16467 &  n_32078;
assign n_32080 = ~n_16461 &  n_32079;
assign n_32081 = ~n_16455 &  n_32080;
assign n_32082 = ~n_16449 &  n_32081;
assign n_32083 = ~n_16443 &  n_32082;
assign n_32084 = ~n_16437 &  n_32083;
assign n_32085 = ~n_16431 &  n_32084;
assign n_32086 = ~n_16425 &  n_32085;
assign n_32087 = ~n_16419 &  n_32086;
assign n_32088 = ~n_16413 &  n_32087;
assign n_32089 = ~n_16407 &  n_32088;
assign n_32090 = ~n_16401 &  n_32089;
assign n_32091 = ~n_16395 &  n_32090;
assign n_32092 = ~n_16389 &  n_32091;
assign n_32093 = ~n_16383 &  n_32092;
assign n_32094 = ~n_16377 &  n_32093;
assign n_32095 = ~n_16371 &  n_32094;
assign n_32096 = ~n_16365 &  n_32095;
assign n_32097 = ~n_16359 &  n_32096;
assign n_32098 = ~n_16353 &  n_32097;
assign n_32099 = ~n_16347 &  n_32098;
assign n_32100 = ~n_16341 &  n_32099;
assign n_32101 = ~n_16333 &  n_32100;
assign n_32102 = ~n_16327 &  n_32101;
assign n_32103 = ~n_16321 &  n_32102;
assign n_32104 = ~n_16315 &  n_32103;
assign n_32105 = ~n_16309 &  n_32104;
assign n_32106 = ~n_16303 &  n_32105;
assign n_32107 = ~n_16297 &  n_32106;
assign n_32108 = ~n_16291 &  n_32107;
assign n_32109 = ~n_16285 &  n_32108;
assign n_32110 = ~n_16279 &  n_32109;
assign n_32111 = ~n_16273 &  n_32110;
assign n_32112 = ~n_16267 &  n_32111;
assign n_32113 = ~n_16261 &  n_32112;
assign n_32114 = ~n_16255 &  n_32113;
assign n_32115 = ~n_16249 &  n_32114;
assign n_32116 = ~n_16243 &  n_32115;
assign n_32117 = ~n_16237 &  n_32116;
assign n_32118 = ~n_16231 &  n_32117;
assign n_32119 = ~n_16225 &  n_32118;
assign n_32120 = ~n_16219 &  n_32119;
assign n_32121 = ~n_16213 &  n_32120;
assign n_32122 = ~n_16207 &  n_32121;
assign n_32123 = ~n_16201 &  n_32122;
assign n_32124 = ~n_16195 &  n_32123;
assign n_32125 = ~n_16189 &  n_32124;
assign n_32126 = ~n_16183 &  n_32125;
assign n_32127 = ~n_16177 &  n_32126;
assign n_32128 = ~n_16171 &  n_32127;
assign n_32129 = ~n_16165 &  n_32128;
assign n_32130 = ~n_16159 &  n_32129;
assign n_32131 = ~n_16153 &  n_32130;
assign n_32132 = ~n_16147 &  n_32131;
assign n_32133 = ~n_16140 &  n_32132;
assign n_32134 = ~n_16134 &  n_32133;
assign n_32135 = ~n_16128 &  n_32134;
assign n_32136 = ~n_16122 &  n_32135;
assign n_32137 = ~n_16116 &  n_32136;
assign n_32138 = ~n_16110 &  n_32137;
assign n_32139 = ~n_16104 &  n_32138;
assign n_32140 = ~n_16098 &  n_32139;
assign n_32141 = ~n_16092 &  n_32140;
assign n_32142 = ~n_16086 &  n_32141;
assign n_32143 = ~n_16080 &  n_32142;
assign n_32144 = ~n_16074 &  n_32143;
assign n_32145 = ~n_16068 &  n_32144;
assign n_32146 = ~n_16062 &  n_32145;
assign n_32147 = ~n_16056 &  n_32146;
assign n_32148 = ~n_16050 &  n_32147;
assign n_32149 = ~n_16044 &  n_32148;
assign n_32150 = ~n_16038 &  n_32149;
assign n_32151 = ~n_16032 &  n_32150;
assign n_32152 = ~n_16026 &  n_32151;
assign n_32153 = ~n_16020 &  n_32152;
assign n_32154 = ~n_16014 &  n_32153;
assign n_32155 = ~n_16008 &  n_32154;
assign n_32156 = ~n_16002 &  n_32155;
assign n_32157 = ~n_15996 &  n_32156;
assign n_32158 = ~n_15990 &  n_32157;
assign n_32159 = ~n_15984 &  n_32158;
assign n_32160 = ~n_15978 &  n_32159;
assign n_32161 = ~n_15972 &  n_32160;
assign n_32162 = ~n_15966 &  n_32161;
assign n_32163 = ~n_15960 &  n_32162;
assign n_32164 = ~n_15954 &  n_32163;
assign n_32165 = ~n_15947 &  n_32164;
assign n_32166 = ~n_15941 &  n_32165;
assign n_32167 = ~n_15935 &  n_32166;
assign n_32168 = ~n_15929 &  n_32167;
assign n_32169 = ~n_15923 &  n_32168;
assign n_32170 = ~n_15917 &  n_32169;
assign n_32171 = ~n_15911 &  n_32170;
assign n_32172 = ~n_15905 &  n_32171;
assign n_32173 = ~n_15899 &  n_32172;
assign n_32174 = ~n_15893 &  n_32173;
assign n_32175 = ~n_15887 &  n_32174;
assign n_32176 = ~n_15881 &  n_32175;
assign n_32177 = ~n_15875 &  n_32176;
assign n_32178 = ~n_15869 &  n_32177;
assign n_32179 = ~n_15863 &  n_32178;
assign n_32180 = ~n_15857 &  n_32179;
assign n_32181 = ~n_15851 &  n_32180;
assign n_32182 = ~n_15845 &  n_32181;
assign n_32183 = ~n_15839 &  n_32182;
assign n_32184 = ~n_15833 &  n_32183;
assign n_32185 = ~n_15827 &  n_32184;
assign n_32186 = ~n_15821 &  n_32185;
assign n_32187 = ~n_15815 &  n_32186;
assign n_32188 = ~n_15809 &  n_32187;
assign n_32189 = ~n_15803 &  n_32188;
assign n_32190 = ~n_15797 &  n_32189;
assign n_32191 = ~n_15791 &  n_32190;
assign n_32192 = ~n_15785 &  n_32191;
assign n_32193 = ~n_15779 &  n_32192;
assign n_32194 = ~n_15773 &  n_32193;
assign n_32195 = ~n_15767 &  n_32194;
assign n_32196 = ~n_15761 &  n_32195;
assign n_32197 = ~n_15754 &  n_32196;
assign n_32198 = ~n_15726 &  n_32197;
assign n_32199 = ~n_15696 &  n_32198;
assign n_32200 = ~n_15666 &  n_32199;
assign n_32201 = ~n_15636 &  n_32200;
assign n_32202 = ~n_15606 &  n_32201;
assign n_32203 = ~n_15576 &  n_32202;
assign n_32204 = ~n_15546 &  n_32203;
assign n_32205 = ~n_15516 &  n_32204;
assign n_32206 = ~n_15486 &  n_32205;
assign n_32207 = ~n_15456 &  n_32206;
assign n_32208 = ~n_15426 &  n_32207;
assign n_32209 = ~n_15396 &  n_32208;
assign n_32210 = ~n_15366 &  n_32209;
assign n_32211 = ~n_15336 &  n_32210;
assign n_32212 = ~n_15306 &  n_32211;
assign n_32213 = ~n_15276 &  n_32212;
assign n_32214 = ~n_15246 &  n_32213;
assign n_32215 = ~n_15216 &  n_32214;
assign n_32216 = ~n_15186 &  n_32215;
assign n_32217 = ~n_15156 &  n_32216;
assign n_32218 = ~n_15126 &  n_32217;
assign n_32219 = ~n_15096 &  n_32218;
assign n_32220 = ~n_15066 &  n_32219;
assign n_32221 = ~n_15036 &  n_32220;
assign n_32222 = ~n_15006 &  n_32221;
assign n_32223 = ~n_14976 &  n_32222;
assign n_32224 = ~n_14946 &  n_32223;
assign n_32225 = ~n_14916 &  n_32224;
assign n_32226 = ~n_14886 &  n_32225;
assign n_32227 = ~n_14852 &  n_32226;
assign n_32228 = ~n_14826 &  n_32227;
assign n_32229 = ~n_14806 &  n_32228;
assign n_32230 = ~n_14778 &  n_32229;
assign n_32231 = ~n_14748 &  n_32230;
assign n_32232 = ~n_14718 &  n_32231;
assign n_32233 = ~n_14688 &  n_32232;
assign n_32234 = ~n_14658 &  n_32233;
assign n_32235 = ~n_14628 &  n_32234;
assign n_32236 = ~n_14598 &  n_32235;
assign n_32237 = ~n_14568 &  n_32236;
assign n_32238 = ~n_14538 &  n_32237;
assign n_32239 = ~n_14508 &  n_32238;
assign n_32240 = ~n_14478 &  n_32239;
assign n_32241 = ~n_14448 &  n_32240;
assign n_32242 = ~n_14418 &  n_32241;
assign n_32243 = ~n_14388 &  n_32242;
assign n_32244 = ~n_14358 &  n_32243;
assign n_32245 = ~n_14328 &  n_32244;
assign n_32246 = ~n_14298 &  n_32245;
assign n_32247 = ~n_14268 &  n_32246;
assign n_32248 = ~n_14238 &  n_32247;
assign n_32249 = ~n_14208 &  n_32248;
assign n_32250 = ~n_14178 &  n_32249;
assign n_32251 = ~n_14148 &  n_32250;
assign n_32252 = ~n_14118 &  n_32251;
assign n_32253 = ~n_14088 &  n_32252;
assign n_32254 = ~n_14058 &  n_32253;
assign n_32255 = ~n_14028 &  n_32254;
assign n_32256 = ~n_13998 &  n_32255;
assign n_32257 = ~n_13968 &  n_32256;
assign n_32258 = ~n_13938 &  n_32257;
assign n_32259 = ~n_13904 &  n_32258;
assign n_32260 = ~n_13878 &  n_32259;
assign n_32261 = ~n_13859 &  n_32260;
assign n_32262 = ~n_13853 &  n_32261;
assign n_32263 = ~n_13847 &  n_32262;
assign n_32264 = ~n_13841 &  n_32263;
assign n_32265 = ~n_13835 &  n_32264;
assign n_32266 = ~n_13829 &  n_32265;
assign n_32267 = ~n_13823 &  n_32266;
assign n_32268 = ~n_13817 &  n_32267;
assign n_32269 = ~n_13811 &  n_32268;
assign n_32270 = ~n_13805 &  n_32269;
assign n_32271 = ~n_13799 &  n_32270;
assign n_32272 = ~n_13793 &  n_32271;
assign n_32273 = ~n_13787 &  n_32272;
assign n_32274 = ~n_13781 &  n_32273;
assign n_32275 = ~n_13775 &  n_32274;
assign n_32276 = ~n_13769 &  n_32275;
assign n_32277 = ~n_13763 &  n_32276;
assign n_32278 = ~n_13757 &  n_32277;
assign n_32279 = ~n_13751 &  n_32278;
assign n_32280 = ~n_13745 &  n_32279;
assign n_32281 = ~n_13739 &  n_32280;
assign n_32282 = ~n_13733 &  n_32281;
assign n_32283 = ~n_13727 &  n_32282;
assign n_32284 = ~n_13721 &  n_32283;
assign n_32285 = ~n_13715 &  n_32284;
assign n_32286 = ~n_13709 &  n_32285;
assign n_32287 = ~n_13703 &  n_32286;
assign n_32288 = ~n_13697 &  n_32287;
assign n_32289 = ~n_13691 &  n_32288;
assign n_32290 = ~n_13685 &  n_32289;
assign n_32291 = ~n_13679 &  n_32290;
assign n_32292 = ~n_13673 &  n_32291;
assign n_32293 = ~n_13666 &  n_32292;
assign n_32294 = ~n_13660 &  n_32293;
assign n_32295 = ~n_13654 &  n_32294;
assign n_32296 = ~n_13648 &  n_32295;
assign n_32297 = ~n_13642 &  n_32296;
assign n_32298 = ~n_13636 &  n_32297;
assign n_32299 = ~n_13630 &  n_32298;
assign n_32300 = ~n_13624 &  n_32299;
assign n_32301 = ~n_13618 &  n_32300;
assign n_32302 = ~n_13612 &  n_32301;
assign n_32303 = ~n_13606 &  n_32302;
assign n_32304 = ~n_13600 &  n_32303;
assign n_32305 = ~n_13594 &  n_32304;
assign n_32306 = ~n_13588 &  n_32305;
assign n_32307 = ~n_13582 &  n_32306;
assign n_32308 = ~n_13576 &  n_32307;
assign n_32309 = ~n_13570 &  n_32308;
assign n_32310 = ~n_13564 &  n_32309;
assign n_32311 = ~n_13558 &  n_32310;
assign n_32312 = ~n_13552 &  n_32311;
assign n_32313 = ~n_13546 &  n_32312;
assign n_32314 = ~n_13540 &  n_32313;
assign n_32315 = ~n_13534 &  n_32314;
assign n_32316 = ~n_13528 &  n_32315;
assign n_32317 = ~n_13522 &  n_32316;
assign n_32318 = ~n_13516 &  n_32317;
assign n_32319 = ~n_13510 &  n_32318;
assign n_32320 = ~n_13504 &  n_32319;
assign n_32321 = ~n_13498 &  n_32320;
assign n_32322 = ~n_13492 &  n_32321;
assign n_32323 = ~n_13486 &  n_32322;
assign n_32324 = ~n_13480 &  n_32323;
assign n_32325 = ~n_13472 &  n_32324;
assign n_32326 = ~n_13458 &  n_32325;
assign n_32327 = ~n_13444 &  n_32326;
assign n_32328 = ~n_13430 &  n_32327;
assign n_32329 = ~n_13416 &  n_32328;
assign n_32330 = ~n_13402 &  n_32329;
assign n_32331 = ~n_13388 &  n_32330;
assign n_32332 = ~n_13374 &  n_32331;
assign n_32333 = ~n_13360 &  n_32332;
assign n_32334 = ~n_13346 &  n_32333;
assign n_32335 = ~n_13332 &  n_32334;
assign n_32336 = ~n_13318 &  n_32335;
assign n_32337 = ~n_13304 &  n_32336;
assign n_32338 = ~n_13290 &  n_32337;
assign n_32339 = ~n_13276 &  n_32338;
assign n_32340 = ~n_13262 &  n_32339;
assign n_32341 = ~n_13248 &  n_32340;
assign n_32342 = ~n_13234 &  n_32341;
assign n_32343 = ~n_13220 &  n_32342;
assign n_32344 = ~n_13206 &  n_32343;
assign n_32345 = ~n_13192 &  n_32344;
assign n_32346 = ~n_13178 &  n_32345;
assign n_32347 = ~n_13164 &  n_32346;
assign n_32348 = ~n_13150 &  n_32347;
assign n_32349 = ~n_13136 &  n_32348;
assign n_32350 = ~n_13122 &  n_32349;
assign n_32351 = ~n_13108 &  n_32350;
assign n_32352 = ~n_13094 &  n_32351;
assign n_32353 = ~n_13080 &  n_32352;
assign n_32354 = ~n_13066 &  n_32353;
assign n_32355 = ~n_13052 &  n_32354;
assign n_32356 = ~n_13038 &  n_32355;
assign n_32357 = ~n_13001 &  n_32356;
assign n_32358 = ~n_12995 &  n_32357;
assign n_32359 = ~n_12989 &  n_32358;
assign n_32360 = ~n_12983 &  n_32359;
assign n_32361 = ~n_12977 &  n_32360;
assign n_32362 = ~n_12971 &  n_32361;
assign n_32363 = ~n_12965 &  n_32362;
assign n_32364 = ~n_12959 &  n_32363;
assign n_32365 = ~n_12953 &  n_32364;
assign n_32366 = ~n_12947 &  n_32365;
assign n_32367 = ~n_12941 &  n_32366;
assign n_32368 = ~n_12935 &  n_32367;
assign n_32369 = ~n_12929 &  n_32368;
assign n_32370 = ~n_12923 &  n_32369;
assign n_32371 = ~n_12917 &  n_32370;
assign n_32372 = ~n_12911 &  n_32371;
assign n_32373 = ~n_12905 &  n_32372;
assign n_32374 = ~n_12899 &  n_32373;
assign n_32375 = ~n_12893 &  n_32374;
assign n_32376 = ~n_12887 &  n_32375;
assign n_32377 = ~n_12881 &  n_32376;
assign n_32378 = ~n_12875 &  n_32377;
assign n_32379 = ~n_12869 &  n_32378;
assign n_32380 = ~n_12863 &  n_32379;
assign n_32381 = ~n_12857 &  n_32380;
assign n_32382 = ~n_12851 &  n_32381;
assign n_32383 = ~n_12845 &  n_32382;
assign n_32384 = ~n_12839 &  n_32383;
assign n_32385 = ~n_12833 &  n_32384;
assign n_32386 = ~n_12827 &  n_32385;
assign n_32387 = ~n_12821 &  n_32386;
assign n_32388 = ~n_12815 &  n_32387;
assign n_32389 = ~n_12808 &  n_32388;
assign n_32390 = ~n_12802 &  n_32389;
assign n_32391 = ~n_12796 &  n_32390;
assign n_32392 = ~n_12790 &  n_32391;
assign n_32393 = ~n_12784 &  n_32392;
assign n_32394 = ~n_12778 &  n_32393;
assign n_32395 = ~n_12772 &  n_32394;
assign n_32396 = ~n_12766 &  n_32395;
assign n_32397 = ~n_12760 &  n_32396;
assign n_32398 = ~n_12754 &  n_32397;
assign n_32399 = ~n_12748 &  n_32398;
assign n_32400 = ~n_12742 &  n_32399;
assign n_32401 = ~n_12736 &  n_32400;
assign n_32402 = ~n_12730 &  n_32401;
assign n_32403 = ~n_12724 &  n_32402;
assign n_32404 = ~n_12718 &  n_32403;
assign n_32405 = ~n_12712 &  n_32404;
assign n_32406 = ~n_12706 &  n_32405;
assign n_32407 = ~n_12700 &  n_32406;
assign n_32408 = ~n_12694 &  n_32407;
assign n_32409 = ~n_12688 &  n_32408;
assign n_32410 = ~n_12682 &  n_32409;
assign n_32411 = ~n_12676 &  n_32410;
assign n_32412 = ~n_12670 &  n_32411;
assign n_32413 = ~n_12664 &  n_32412;
assign n_32414 = ~n_12658 &  n_32413;
assign n_32415 = ~n_12652 &  n_32414;
assign n_32416 = ~n_12646 &  n_32415;
assign n_32417 = ~n_12640 &  n_32416;
assign n_32418 = ~n_12634 &  n_32417;
assign n_32419 = ~n_12628 &  n_32418;
assign n_32420 = ~n_12622 &  n_32419;
assign n_32421 = ~n_12613 &  n_32420;
assign n_32422 = ~n_12607 &  n_32421;
assign n_32423 = ~n_12601 &  n_32422;
assign n_32424 = ~n_12595 &  n_32423;
assign n_32425 = ~n_12589 &  n_32424;
assign n_32426 = ~n_12583 &  n_32425;
assign n_32427 = ~n_12577 &  n_32426;
assign n_32428 = ~n_12571 &  n_32427;
assign n_32429 = ~n_12565 &  n_32428;
assign n_32430 = ~n_12559 &  n_32429;
assign n_32431 = ~n_12553 &  n_32430;
assign n_32432 = ~n_12547 &  n_32431;
assign n_32433 = ~n_12541 &  n_32432;
assign n_32434 = ~n_12535 &  n_32433;
assign n_32435 = ~n_12529 &  n_32434;
assign n_32436 = ~n_12523 &  n_32435;
assign n_32437 = ~n_12517 &  n_32436;
assign n_32438 = ~n_12511 &  n_32437;
assign n_32439 = ~n_12505 &  n_32438;
assign n_32440 = ~n_12499 &  n_32439;
assign n_32441 = ~n_12493 &  n_32440;
assign n_32442 = ~n_12487 &  n_32441;
assign n_32443 = ~n_12481 &  n_32442;
assign n_32444 = ~n_12475 &  n_32443;
assign n_32445 = ~n_12469 &  n_32444;
assign n_32446 = ~n_12463 &  n_32445;
assign n_32447 = ~n_12457 &  n_32446;
assign n_32448 = ~n_12451 &  n_32447;
assign n_32449 = ~n_12445 &  n_32448;
assign n_32450 = ~n_12439 &  n_32449;
assign n_32451 = ~n_12433 &  n_32450;
assign n_32452 = ~n_12427 &  n_32451;
assign n_32453 = ~n_12419 &  n_32452;
assign n_32454 = ~n_12413 &  n_32453;
assign n_32455 = ~n_12407 &  n_32454;
assign n_32456 = ~n_12401 &  n_32455;
assign n_32457 = ~n_12395 &  n_32456;
assign n_32458 = ~n_12389 &  n_32457;
assign n_32459 = ~n_12383 &  n_32458;
assign n_32460 = ~n_12377 &  n_32459;
assign n_32461 = ~n_12371 &  n_32460;
assign n_32462 = ~n_12365 &  n_32461;
assign n_32463 = ~n_12359 &  n_32462;
assign n_32464 = ~n_12353 &  n_32463;
assign n_32465 = ~n_12347 &  n_32464;
assign n_32466 = ~n_12341 &  n_32465;
assign n_32467 = ~n_12335 &  n_32466;
assign n_32468 = ~n_12329 &  n_32467;
assign n_32469 = ~n_12323 &  n_32468;
assign n_32470 = ~n_12317 &  n_32469;
assign n_32471 = ~n_12311 &  n_32470;
assign n_32472 = ~n_12305 &  n_32471;
assign n_32473 = ~n_12299 &  n_32472;
assign n_32474 = ~n_12293 &  n_32473;
assign n_32475 = ~n_12287 &  n_32474;
assign n_32476 = ~n_12281 &  n_32475;
assign n_32477 = ~n_12275 &  n_32476;
assign n_32478 = ~n_12269 &  n_32477;
assign n_32479 = ~n_12263 &  n_32478;
assign n_32480 = ~n_12257 &  n_32479;
assign n_32481 = ~n_12251 &  n_32480;
assign n_32482 = ~n_12245 &  n_32481;
assign n_32483 = ~n_12239 &  n_32482;
assign n_32484 = ~n_12233 &  n_32483;
assign n_32485 = ~n_12225 &  n_32484;
assign n_32486 = ~n_12219 &  n_32485;
assign n_32487 = ~n_12213 &  n_32486;
assign n_32488 = ~n_12207 &  n_32487;
assign n_32489 = ~n_12201 &  n_32488;
assign n_32490 = ~n_12195 &  n_32489;
assign n_32491 = ~n_12189 &  n_32490;
assign n_32492 = ~n_12183 &  n_32491;
assign n_32493 = ~n_12177 &  n_32492;
assign n_32494 = ~n_12171 &  n_32493;
assign n_32495 = ~n_12165 &  n_32494;
assign n_32496 = ~n_12159 &  n_32495;
assign n_32497 = ~n_12153 &  n_32496;
assign n_32498 = ~n_12147 &  n_32497;
assign n_32499 = ~n_12141 &  n_32498;
assign n_32500 = ~n_12135 &  n_32499;
assign n_32501 = ~n_12129 &  n_32500;
assign n_32502 = ~n_12123 &  n_32501;
assign n_32503 = ~n_12117 &  n_32502;
assign n_32504 = ~n_12111 &  n_32503;
assign n_32505 = ~n_12105 &  n_32504;
assign n_32506 = ~n_12099 &  n_32505;
assign n_32507 = ~n_12093 &  n_32506;
assign n_32508 = ~n_12087 &  n_32507;
assign n_32509 = ~n_12081 &  n_32508;
assign n_32510 = ~n_12075 &  n_32509;
assign n_32511 = ~n_12069 &  n_32510;
assign n_32512 = ~n_12063 &  n_32511;
assign n_32513 = ~n_12057 &  n_32512;
assign n_32514 = ~n_12051 &  n_32513;
assign n_32515 = ~n_12045 &  n_32514;
assign n_32516 = ~n_12039 &  n_32515;
assign n_32517 = ~n_12031 &  n_32516;
assign n_32518 = ~n_11986 &  n_32517;
assign n_32519 = ~n_11938 &  n_32518;
assign n_32520 = ~n_11890 &  n_32519;
assign n_32521 = ~n_11842 &  n_32520;
assign n_32522 = ~n_11794 &  n_32521;
assign n_32523 = ~n_11746 &  n_32522;
assign n_32524 = ~n_11698 &  n_32523;
assign n_32525 = ~n_11650 &  n_32524;
assign n_32526 = ~n_11602 &  n_32525;
assign n_32527 = ~n_11554 &  n_32526;
assign n_32528 = ~n_11506 &  n_32527;
assign n_32529 = ~n_11458 &  n_32528;
assign n_32530 = ~n_11410 &  n_32529;
assign n_32531 = ~n_11362 &  n_32530;
assign n_32532 = ~n_11314 &  n_32531;
assign n_32533 = ~n_11266 &  n_32532;
assign n_32534 = ~n_11218 &  n_32533;
assign n_32535 = ~n_11170 &  n_32534;
assign n_32536 = ~n_11122 &  n_32535;
assign n_32537 = ~n_11074 &  n_32536;
assign n_32538 = ~n_11026 &  n_32537;
assign n_32539 = ~n_10978 &  n_32538;
assign n_32540 = ~n_10930 &  n_32539;
assign n_32541 = ~n_10882 &  n_32540;
assign n_32542 = ~n_10834 &  n_32541;
assign n_32543 = ~n_10786 &  n_32542;
assign n_32544 = ~n_10738 &  n_32543;
assign n_32545 = ~n_10690 &  n_32544;
assign n_32546 = ~n_10642 &  n_32545;
assign n_32547 = ~n_10588 &  n_32546;
assign n_32548 = ~n_10546 &  n_32547;
assign n_32549 = ~n_10514 &  n_32548;
assign n_32550 = ~n_10508 &  n_32549;
assign n_32551 = ~n_10502 &  n_32550;
assign n_32552 = ~n_10496 &  n_32551;
assign n_32553 = ~n_10490 &  n_32552;
assign n_32554 = ~n_10484 &  n_32553;
assign n_32555 = ~n_10478 &  n_32554;
assign n_32556 = ~n_10472 &  n_32555;
assign n_32557 = ~n_10466 &  n_32556;
assign n_32558 = ~n_10460 &  n_32557;
assign n_32559 = ~n_10454 &  n_32558;
assign n_32560 = ~n_10448 &  n_32559;
assign n_32561 = ~n_10442 &  n_32560;
assign n_32562 = ~n_10436 &  n_32561;
assign n_32563 = ~n_10430 &  n_32562;
assign n_32564 = ~n_10424 &  n_32563;
assign n_32565 = ~n_10418 &  n_32564;
assign n_32566 = ~n_10412 &  n_32565;
assign n_32567 = ~n_10406 &  n_32566;
assign n_32568 = ~n_10400 &  n_32567;
assign n_32569 = ~n_10394 &  n_32568;
assign n_32570 = ~n_10388 &  n_32569;
assign n_32571 = ~n_10382 &  n_32570;
assign n_32572 = ~n_10376 &  n_32571;
assign n_32573 = ~n_10370 &  n_32572;
assign n_32574 = ~n_10364 &  n_32573;
assign n_32575 = ~n_10358 &  n_32574;
assign n_32576 = ~n_10352 &  n_32575;
assign n_32577 = ~n_10346 &  n_32576;
assign n_32578 = ~n_10340 &  n_32577;
assign n_32579 = ~n_10334 &  n_32578;
assign n_32580 = ~n_10328 &  n_32579;
assign n_32581 = ~n_10317 &  n_32580;
assign n_32582 = ~n_10271 &  n_32581;
assign n_32583 = ~n_10223 &  n_32582;
assign n_32584 = ~n_10175 &  n_32583;
assign n_32585 = ~n_10127 &  n_32584;
assign n_32586 = ~n_10079 &  n_32585;
assign n_32587 = ~n_10031 &  n_32586;
assign n_32588 = ~n_9983 &  n_32587;
assign n_32589 = ~n_9935 &  n_32588;
assign n_32590 = ~n_9887 &  n_32589;
assign n_32591 = ~n_9839 &  n_32590;
assign n_32592 = ~n_9791 &  n_32591;
assign n_32593 = ~n_9743 &  n_32592;
assign n_32594 = ~n_9695 &  n_32593;
assign n_32595 = ~n_9647 &  n_32594;
assign n_32596 = ~n_9599 &  n_32595;
assign n_32597 = ~n_9551 &  n_32596;
assign n_32598 = ~n_9503 &  n_32597;
assign n_32599 = ~n_9455 &  n_32598;
assign n_32600 = ~n_9407 &  n_32599;
assign n_32601 = ~n_9359 &  n_32600;
assign n_32602 = ~n_9311 &  n_32601;
assign n_32603 = ~n_9263 &  n_32602;
assign n_32604 = ~n_9215 &  n_32603;
assign n_32605 = ~n_9167 &  n_32604;
assign n_32606 = ~n_9119 &  n_32605;
assign n_32607 = ~n_9071 &  n_32606;
assign n_32608 = ~n_9023 &  n_32607;
assign n_32609 = ~n_8975 &  n_32608;
assign n_32610 = ~n_8927 &  n_32609;
assign n_32611 = ~n_8874 &  n_32610;
assign n_32612 = ~n_8832 &  n_32611;
assign n_32613 = ~n_8801 &  n_32612;
assign n_32614 = ~n_8796 &  n_32613;
assign n_32615 = ~n_8791 &  n_32614;
assign n_32616 = ~n_8786 &  n_32615;
assign n_32617 = ~n_8781 &  n_32616;
assign n_32618 = ~n_8776 &  n_32617;
assign n_32619 = ~n_8771 &  n_32618;
assign n_32620 = ~n_8766 &  n_32619;
assign n_32621 = ~n_8761 &  n_32620;
assign n_32622 = ~n_8756 &  n_32621;
assign n_32623 = ~n_8751 &  n_32622;
assign n_32624 = ~n_8746 &  n_32623;
assign n_32625 = ~n_8741 &  n_32624;
assign n_32626 = ~n_8736 &  n_32625;
assign n_32627 = ~n_8731 &  n_32626;
assign n_32628 = ~n_8726 &  n_32627;
assign n_32629 = ~n_8721 &  n_32628;
assign n_32630 = ~n_8716 &  n_32629;
assign n_32631 = ~n_8711 &  n_32630;
assign n_32632 = ~n_8706 &  n_32631;
assign n_32633 = ~n_8701 &  n_32632;
assign n_32634 = ~n_8696 &  n_32633;
assign n_32635 = ~n_8691 &  n_32634;
assign n_32636 = ~n_8686 &  n_32635;
assign n_32637 = ~n_8681 &  n_32636;
assign n_32638 = ~n_8676 &  n_32637;
assign n_32639 = ~n_8671 &  n_32638;
assign n_32640 = ~n_8666 &  n_32639;
assign n_32641 = ~n_8661 &  n_32640;
assign n_32642 = ~n_8656 &  n_32641;
assign n_32643 = ~n_8651 &  n_32642;
assign n_32644 = ~n_8646 &  n_32643;
assign n_32645 = ~n_8641 &  n_32644;
assign n_32646 = ~n_8635 &  n_32645;
assign n_32647 = ~n_8629 &  n_32646;
assign n_32648 = ~n_8623 &  n_32647;
assign n_32649 = ~n_8617 &  n_32648;
assign n_32650 = ~n_8611 &  n_32649;
assign n_32651 = ~n_8605 &  n_32650;
assign n_32652 = ~n_8599 &  n_32651;
assign n_32653 = ~n_8593 &  n_32652;
assign n_32654 = ~n_8587 &  n_32653;
assign n_32655 = ~n_8581 &  n_32654;
assign n_32656 = ~n_8575 &  n_32655;
assign n_32657 = ~n_8569 &  n_32656;
assign n_32658 = ~n_8563 &  n_32657;
assign n_32659 = ~n_8557 &  n_32658;
assign n_32660 = ~n_8551 &  n_32659;
assign n_32661 = ~n_8545 &  n_32660;
assign n_32662 = ~n_8539 &  n_32661;
assign n_32663 = ~n_8533 &  n_32662;
assign n_32664 = ~n_8527 &  n_32663;
assign n_32665 = ~n_8521 &  n_32664;
assign n_32666 = ~n_8515 &  n_32665;
assign n_32667 = ~n_8509 &  n_32666;
assign n_32668 = ~n_8503 &  n_32667;
assign n_32669 = ~n_8497 &  n_32668;
assign n_32670 = ~n_8491 &  n_32669;
assign n_32671 = ~n_8485 &  n_32670;
assign n_32672 = ~n_8479 &  n_32671;
assign n_32673 = ~n_8473 &  n_32672;
assign n_32674 = ~n_8467 &  n_32673;
assign n_32675 = ~n_8461 &  n_32674;
assign n_32676 = ~n_8455 &  n_32675;
assign n_32677 = ~n_8448 &  n_32676;
assign n_32678 = ~n_8442 &  n_32677;
assign n_32679 = ~n_8436 &  n_32678;
assign n_32680 = ~n_8430 &  n_32679;
assign n_32681 = ~n_8424 &  n_32680;
assign n_32682 = ~n_8418 &  n_32681;
assign n_32683 = ~n_8412 &  n_32682;
assign n_32684 = ~n_8406 &  n_32683;
assign n_32685 = ~n_8400 &  n_32684;
assign n_32686 = ~n_8394 &  n_32685;
assign n_32687 = ~n_8388 &  n_32686;
assign n_32688 = ~n_8382 &  n_32687;
assign n_32689 = ~n_8376 &  n_32688;
assign n_32690 = ~n_8370 &  n_32689;
assign n_32691 = ~n_8364 &  n_32690;
assign n_32692 = ~n_8358 &  n_32691;
assign n_32693 = ~n_8352 &  n_32692;
assign n_32694 = ~n_8346 &  n_32693;
assign n_32695 = ~n_8340 &  n_32694;
assign n_32696 = ~n_8334 &  n_32695;
assign n_32697 = ~n_8328 &  n_32696;
assign n_32698 = ~n_8322 &  n_32697;
assign n_32699 = ~n_8316 &  n_32698;
assign n_32700 = ~n_8310 &  n_32699;
assign n_32701 = ~n_8304 &  n_32700;
assign n_32702 = ~n_8298 &  n_32701;
assign n_32703 = ~n_8292 &  n_32702;
assign n_32704 = ~n_8286 &  n_32703;
assign n_32705 = ~n_8280 &  n_32704;
assign n_32706 = ~n_8274 &  n_32705;
assign n_32707 = ~n_8268 &  n_32706;
assign n_32708 = ~n_8262 &  n_32707;
assign n_32709 = ~n_8253 &  n_32708;
assign n_32710 = ~n_8247 &  n_32709;
assign n_32711 = ~n_8241 &  n_32710;
assign n_32712 = ~n_8235 &  n_32711;
assign n_32713 = ~n_8229 &  n_32712;
assign n_32714 = ~n_8223 &  n_32713;
assign n_32715 = ~n_8217 &  n_32714;
assign n_32716 = ~n_8211 &  n_32715;
assign n_32717 = ~n_8205 &  n_32716;
assign n_32718 = ~n_8199 &  n_32717;
assign n_32719 = ~n_8193 &  n_32718;
assign n_32720 = ~n_8187 &  n_32719;
assign n_32721 = ~n_8181 &  n_32720;
assign n_32722 = ~n_8175 &  n_32721;
assign n_32723 = ~n_8169 &  n_32722;
assign n_32724 = ~n_8163 &  n_32723;
assign n_32725 = ~n_8157 &  n_32724;
assign n_32726 = ~n_8151 &  n_32725;
assign n_32727 = ~n_8145 &  n_32726;
assign n_32728 = ~n_8139 &  n_32727;
assign n_32729 = ~n_8133 &  n_32728;
assign n_32730 = ~n_8127 &  n_32729;
assign n_32731 = ~n_8121 &  n_32730;
assign n_32732 = ~n_8115 &  n_32731;
assign n_32733 = ~n_8109 &  n_32732;
assign n_32734 = ~n_8103 &  n_32733;
assign n_32735 = ~n_8097 &  n_32734;
assign n_32736 = ~n_8091 &  n_32735;
assign n_32737 = ~n_8085 &  n_32736;
assign n_32738 = ~n_8079 &  n_32737;
assign n_32739 = ~n_8073 &  n_32738;
assign n_32740 = ~n_8067 &  n_32739;
assign n_32741 = ~n_8058 &  n_32740;
assign n_32742 = ~n_8052 &  n_32741;
assign n_32743 = ~n_8046 &  n_32742;
assign n_32744 = ~n_8040 &  n_32743;
assign n_32745 = ~n_8034 &  n_32744;
assign n_32746 = ~n_8028 &  n_32745;
assign n_32747 = ~n_8022 &  n_32746;
assign n_32748 = ~n_8016 &  n_32747;
assign n_32749 = ~n_8010 &  n_32748;
assign n_32750 = ~n_8004 &  n_32749;
assign n_32751 = ~n_7998 &  n_32750;
assign n_32752 = ~n_7992 &  n_32751;
assign n_32753 = ~n_7986 &  n_32752;
assign n_32754 = ~n_7980 &  n_32753;
assign n_32755 = ~n_7974 &  n_32754;
assign n_32756 = ~n_7968 &  n_32755;
assign n_32757 = ~n_7962 &  n_32756;
assign n_32758 = ~n_7956 &  n_32757;
assign n_32759 = ~n_7950 &  n_32758;
assign n_32760 = ~n_7944 &  n_32759;
assign n_32761 = ~n_7938 &  n_32760;
assign n_32762 = ~n_7932 &  n_32761;
assign n_32763 = ~n_7926 &  n_32762;
assign n_32764 = ~n_7920 &  n_32763;
assign n_32765 = ~n_7914 &  n_32764;
assign n_32766 = ~n_7908 &  n_32765;
assign n_32767 = ~n_7902 &  n_32766;
assign n_32768 = ~n_7896 &  n_32767;
assign n_32769 = ~n_7890 &  n_32768;
assign n_32770 = ~n_7884 &  n_32769;
assign n_32771 = ~n_7878 &  n_32770;
assign n_32772 = ~n_7872 &  n_32771;
assign n_32773 = ~n_7864 &  n_32772;
assign n_32774 = ~n_7858 &  n_32773;
assign n_32775 = ~n_7852 &  n_32774;
assign n_32776 = ~n_7846 &  n_32775;
assign n_32777 = ~n_7840 &  n_32776;
assign n_32778 = ~n_7834 &  n_32777;
assign n_32779 = ~n_7828 &  n_32778;
assign n_32780 = ~n_7822 &  n_32779;
assign n_32781 = ~n_7816 &  n_32780;
assign n_32782 = ~n_7810 &  n_32781;
assign n_32783 = ~n_7804 &  n_32782;
assign n_32784 = ~n_7798 &  n_32783;
assign n_32785 = ~n_7792 &  n_32784;
assign n_32786 = ~n_7786 &  n_32785;
assign n_32787 = ~n_7780 &  n_32786;
assign n_32788 = ~n_7774 &  n_32787;
assign n_32789 = ~n_7768 &  n_32788;
assign n_32790 = ~n_7762 &  n_32789;
assign n_32791 = ~n_7756 &  n_32790;
assign n_32792 = ~n_7750 &  n_32791;
assign n_32793 = ~n_7744 &  n_32792;
assign n_32794 = ~n_7738 &  n_32793;
assign n_32795 = ~n_7732 &  n_32794;
assign n_32796 = ~n_7726 &  n_32795;
assign n_32797 = ~n_7720 &  n_32796;
assign n_32798 = ~n_7714 &  n_32797;
assign n_32799 = ~n_7708 &  n_32798;
assign n_32800 = ~n_7702 &  n_32799;
assign n_32801 = ~n_7696 &  n_32800;
assign n_32802 = ~n_7690 &  n_32801;
assign n_32803 = ~n_7684 &  n_32802;
assign n_32804 = ~n_7678 &  n_32803;
assign n_32805 = ~n_7671 &  n_32804;
assign n_32806 = ~n_7665 &  n_32805;
assign n_32807 = ~n_7659 &  n_32806;
assign n_32808 = ~n_7653 &  n_32807;
assign n_32809 = ~n_7647 &  n_32808;
assign n_32810 = ~n_7641 &  n_32809;
assign n_32811 = ~n_7635 &  n_32810;
assign n_32812 = ~n_7629 &  n_32811;
assign n_32813 = ~n_7623 &  n_32812;
assign n_32814 = ~n_7617 &  n_32813;
assign n_32815 = ~n_7611 &  n_32814;
assign n_32816 = ~n_7605 &  n_32815;
assign n_32817 = ~n_7599 &  n_32816;
assign n_32818 = ~n_7593 &  n_32817;
assign n_32819 = ~n_7587 &  n_32818;
assign n_32820 = ~n_7581 &  n_32819;
assign n_32821 = ~n_7575 &  n_32820;
assign n_32822 = ~n_7569 &  n_32821;
assign n_32823 = ~n_7563 &  n_32822;
assign n_32824 = ~n_7557 &  n_32823;
assign n_32825 = ~n_7551 &  n_32824;
assign n_32826 = ~n_7545 &  n_32825;
assign n_32827 = ~n_7539 &  n_32826;
assign n_32828 = ~n_7533 &  n_32827;
assign n_32829 = ~n_7527 &  n_32828;
assign n_32830 = ~n_7521 &  n_32829;
assign n_32831 = ~n_7515 &  n_32830;
assign n_32832 = ~n_7509 &  n_32831;
assign n_32833 = ~n_7503 &  n_32832;
assign n_32834 = ~n_7497 &  n_32833;
assign n_32835 = ~n_7491 &  n_32834;
assign n_32836 = ~n_7485 &  n_32835;
assign n_32837 = ~n_7478 &  n_32836;
assign n_32838 = ~n_7450 &  n_32837;
assign n_32839 = ~n_7420 &  n_32838;
assign n_32840 = ~n_7390 &  n_32839;
assign n_32841 = ~n_7360 &  n_32840;
assign n_32842 = ~n_7330 &  n_32841;
assign n_32843 = ~n_7300 &  n_32842;
assign n_32844 = ~n_7270 &  n_32843;
assign n_32845 = ~n_7240 &  n_32844;
assign n_32846 = ~n_7210 &  n_32845;
assign n_32847 = ~n_7180 &  n_32846;
assign n_32848 = ~n_7150 &  n_32847;
assign n_32849 = ~n_7120 &  n_32848;
assign n_32850 = ~n_7090 &  n_32849;
assign n_32851 = ~n_7060 &  n_32850;
assign n_32852 = ~n_7030 &  n_32851;
assign n_32853 = ~n_7000 &  n_32852;
assign n_32854 = ~n_6970 &  n_32853;
assign n_32855 = ~n_6940 &  n_32854;
assign n_32856 = ~n_6910 &  n_32855;
assign n_32857 = ~n_6880 &  n_32856;
assign n_32858 = ~n_6850 &  n_32857;
assign n_32859 = ~n_6820 &  n_32858;
assign n_32860 = ~n_6790 &  n_32859;
assign n_32861 = ~n_6760 &  n_32860;
assign n_32862 = ~n_6730 &  n_32861;
assign n_32863 = ~n_6700 &  n_32862;
assign n_32864 = ~n_6670 &  n_32863;
assign n_32865 = ~n_6640 &  n_32864;
assign n_32866 = ~n_6610 &  n_32865;
assign n_32867 = ~n_6576 &  n_32866;
assign n_32868 = ~n_6550 &  n_32867;
assign n_32869 = ~n_6526 &  n_32868;
assign n_32870 = ~n_6520 &  n_32869;
assign n_32871 = ~n_6514 &  n_32870;
assign n_32872 = ~n_6508 &  n_32871;
assign n_32873 = ~n_6502 &  n_32872;
assign n_32874 = ~n_6496 &  n_32873;
assign n_32875 = ~n_6490 &  n_32874;
assign n_32876 = ~n_6484 &  n_32875;
assign n_32877 = ~n_6478 &  n_32876;
assign n_32878 = ~n_6472 &  n_32877;
assign n_32879 = ~n_6466 &  n_32878;
assign n_32880 = ~n_6460 &  n_32879;
assign n_32881 = ~n_6454 &  n_32880;
assign n_32882 = ~n_6448 &  n_32881;
assign n_32883 = ~n_6442 &  n_32882;
assign n_32884 = ~n_6436 &  n_32883;
assign n_32885 = ~n_6430 &  n_32884;
assign n_32886 = ~n_6424 &  n_32885;
assign n_32887 = ~n_6418 &  n_32886;
assign n_32888 = ~n_6412 &  n_32887;
assign n_32889 = ~n_6406 &  n_32888;
assign n_32890 = ~n_6400 &  n_32889;
assign n_32891 = ~n_6394 &  n_32890;
assign n_32892 = ~n_6388 &  n_32891;
assign n_32893 = ~n_6382 &  n_32892;
assign n_32894 = ~n_6376 &  n_32893;
assign n_32895 = ~n_6370 &  n_32894;
assign n_32896 = ~n_6364 &  n_32895;
assign n_32897 = ~n_6358 &  n_32896;
assign n_32898 = ~n_6352 &  n_32897;
assign n_32899 = ~n_6346 &  n_32898;
assign n_32900 = ~n_6340 &  n_32899;
assign n_32901 = ~n_6329 &  n_32900;
assign n_32902 = ~n_6323 &  n_32901;
assign n_32903 = ~n_6317 &  n_32902;
assign n_32904 = ~n_6311 &  n_32903;
assign n_32905 = ~n_6305 &  n_32904;
assign n_32906 = ~n_6299 &  n_32905;
assign n_32907 = ~n_6293 &  n_32906;
assign n_32908 = ~n_6287 &  n_32907;
assign n_32909 = ~n_6281 &  n_32908;
assign n_32910 = ~n_6275 &  n_32909;
assign n_32911 = ~n_6269 &  n_32910;
assign n_32912 = ~n_6263 &  n_32911;
assign n_32913 = ~n_6257 &  n_32912;
assign n_32914 = ~n_6251 &  n_32913;
assign n_32915 = ~n_6245 &  n_32914;
assign n_32916 = ~n_6239 &  n_32915;
assign n_32917 = ~n_6233 &  n_32916;
assign n_32918 = ~n_6227 &  n_32917;
assign n_32919 = ~n_6221 &  n_32918;
assign n_32920 = ~n_6215 &  n_32919;
assign n_32921 = ~n_6209 &  n_32920;
assign n_32922 = ~n_6203 &  n_32921;
assign n_32923 = ~n_6197 &  n_32922;
assign n_32924 = ~n_6191 &  n_32923;
assign n_32925 = ~n_6185 &  n_32924;
assign n_32926 = ~n_6179 &  n_32925;
assign n_32927 = ~n_6173 &  n_32926;
assign n_32928 = ~n_6167 &  n_32927;
assign n_32929 = ~n_6161 &  n_32928;
assign n_32930 = ~n_6155 &  n_32929;
assign n_32931 = ~n_6149 &  n_32930;
assign n_32932 = ~n_6143 &  n_32931;
assign n_32933 = ~n_6134 &  n_32932;
assign n_32934 = ~n_6106 &  n_32933;
assign n_32935 = ~n_6076 &  n_32934;
assign n_32936 = ~n_6046 &  n_32935;
assign n_32937 = ~n_6016 &  n_32936;
assign n_32938 = ~n_5986 &  n_32937;
assign n_32939 = ~n_5956 &  n_32938;
assign n_32940 = ~n_5926 &  n_32939;
assign n_32941 = ~n_5896 &  n_32940;
assign n_32942 = ~n_5866 &  n_32941;
assign n_32943 = ~n_5836 &  n_32942;
assign n_32944 = ~n_5806 &  n_32943;
assign n_32945 = ~n_5776 &  n_32944;
assign n_32946 = ~n_5746 &  n_32945;
assign n_32947 = ~n_5716 &  n_32946;
assign n_32948 = ~n_5686 &  n_32947;
assign n_32949 = ~n_5656 &  n_32948;
assign n_32950 = ~n_5626 &  n_32949;
assign n_32951 = ~n_5596 &  n_32950;
assign n_32952 = ~n_5566 &  n_32951;
assign n_32953 = ~n_5536 &  n_32952;
assign n_32954 = ~n_5506 &  n_32953;
assign n_32955 = ~n_5476 &  n_32954;
assign n_32956 = ~n_5446 &  n_32955;
assign n_32957 = ~n_5416 &  n_32956;
assign n_32958 = ~n_5386 &  n_32957;
assign n_32959 = ~n_5356 &  n_32958;
assign n_32960 = ~n_5326 &  n_32959;
assign n_32961 = ~n_5296 &  n_32960;
assign n_32962 = ~n_5266 &  n_32961;
assign n_32963 = ~n_5232 &  n_32962;
assign n_32964 = ~n_5206 &  n_32963;
assign n_32965 = ~n_5186 &  n_32964;
assign n_32966 = ~n_5180 &  n_32965;
assign n_32967 = ~n_5174 &  n_32966;
assign n_32968 = ~n_5168 &  n_32967;
assign n_32969 = ~n_5162 &  n_32968;
assign n_32970 = ~n_5156 &  n_32969;
assign n_32971 = ~n_5150 &  n_32970;
assign n_32972 = ~n_5144 &  n_32971;
assign n_32973 = ~n_5138 &  n_32972;
assign n_32974 = ~n_5132 &  n_32973;
assign n_32975 = ~n_5126 &  n_32974;
assign n_32976 = ~n_5120 &  n_32975;
assign n_32977 = ~n_5114 &  n_32976;
assign n_32978 = ~n_5108 &  n_32977;
assign n_32979 = ~n_5102 &  n_32978;
assign n_32980 = ~n_5096 &  n_32979;
assign n_32981 = ~n_5090 &  n_32980;
assign n_32982 = ~n_5084 &  n_32981;
assign n_32983 = ~n_5078 &  n_32982;
assign n_32984 = ~n_5072 &  n_32983;
assign n_32985 = ~n_5066 &  n_32984;
assign n_32986 = ~n_5060 &  n_32985;
assign n_32987 = ~n_5054 &  n_32986;
assign n_32988 = ~n_5048 &  n_32987;
assign n_32989 = ~n_5042 &  n_32988;
assign n_32990 = ~n_5036 &  n_32989;
assign n_32991 = ~n_5030 &  n_32990;
assign n_32992 = ~n_5024 &  n_32991;
assign n_32993 = ~n_5018 &  n_32992;
assign n_32994 = ~n_5012 &  n_32993;
assign n_32995 = ~n_5006 &  n_32994;
assign n_32996 = ~n_5000 &  n_32995;
assign n_32997 = ~n_4991 &  n_32996;
assign n_32998 = ~n_4986 &  n_32997;
assign n_32999 = ~n_4981 &  n_32998;
assign n_33000 = ~n_4976 &  n_32999;
assign n_33001 = ~n_4971 &  n_33000;
assign n_33002 = ~n_4966 &  n_33001;
assign n_33003 = ~n_4961 &  n_33002;
assign n_33004 = ~n_4956 &  n_33003;
assign n_33005 = ~n_4951 &  n_33004;
assign n_33006 = ~n_4946 &  n_33005;
assign n_33007 = ~n_4941 &  n_33006;
assign n_33008 = ~n_4936 &  n_33007;
assign n_33009 = ~n_4931 &  n_33008;
assign n_33010 = ~n_4926 &  n_33009;
assign n_33011 = ~n_4921 &  n_33010;
assign n_33012 = ~n_4916 &  n_33011;
assign n_33013 = ~n_4911 &  n_33012;
assign n_33014 = ~n_4906 &  n_33013;
assign n_33015 = ~n_4901 &  n_33014;
assign n_33016 = ~n_4896 &  n_33015;
assign n_33017 = ~n_4891 &  n_33016;
assign n_33018 = ~n_4886 &  n_33017;
assign n_33019 = ~n_4881 &  n_33018;
assign n_33020 = ~n_4876 &  n_33019;
assign n_33021 = ~n_4871 &  n_33020;
assign n_33022 = ~n_4866 &  n_33021;
assign n_33023 = ~n_4861 &  n_33022;
assign n_33024 = ~n_4856 &  n_33023;
assign n_33025 = ~n_4851 &  n_33024;
assign n_33026 = ~n_4846 &  n_33025;
assign n_33027 = ~n_4841 &  n_33026;
assign n_33028 = ~n_4836 &  n_33027;
assign n_33029 = ~n_4831 &  n_33028;
assign n_33030 = ~n_4825 &  n_33029;
assign n_33031 = ~n_4819 &  n_33030;
assign n_33032 = ~n_4813 &  n_33031;
assign n_33033 = ~n_4807 &  n_33032;
assign n_33034 = ~n_4801 &  n_33033;
assign n_33035 = ~n_4795 &  n_33034;
assign n_33036 = ~n_4789 &  n_33035;
assign n_33037 = ~n_4783 &  n_33036;
assign n_33038 = ~n_4777 &  n_33037;
assign n_33039 = ~n_4771 &  n_33038;
assign n_33040 = ~n_4765 &  n_33039;
assign n_33041 = ~n_4759 &  n_33040;
assign n_33042 = ~n_4753 &  n_33041;
assign n_33043 = ~n_4747 &  n_33042;
assign n_33044 = ~n_4741 &  n_33043;
assign n_33045 = ~n_4735 &  n_33044;
assign n_33046 = ~n_4729 &  n_33045;
assign n_33047 = ~n_4723 &  n_33046;
assign n_33048 = ~n_4717 &  n_33047;
assign n_33049 = ~n_4711 &  n_33048;
assign n_33050 = ~n_4705 &  n_33049;
assign n_33051 = ~n_4699 &  n_33050;
assign n_33052 = ~n_4693 &  n_33051;
assign n_33053 = ~n_4687 &  n_33052;
assign n_33054 = ~n_4681 &  n_33053;
assign n_33055 = ~n_4675 &  n_33054;
assign n_33056 = ~n_4669 &  n_33055;
assign n_33057 = ~n_4663 &  n_33056;
assign n_33058 = ~n_4657 &  n_33057;
assign n_33059 = ~n_4651 &  n_33058;
assign n_33060 = ~n_4645 &  n_33059;
assign n_33061 = ~n_4638 &  n_33060;
assign n_33062 = ~n_4632 &  n_33061;
assign n_33063 = ~n_4626 &  n_33062;
assign n_33064 = ~n_4620 &  n_33063;
assign n_33065 = ~n_4614 &  n_33064;
assign n_33066 = ~n_4608 &  n_33065;
assign n_33067 = ~n_4602 &  n_33066;
assign n_33068 = ~n_4596 &  n_33067;
assign n_33069 = ~n_4590 &  n_33068;
assign n_33070 = ~n_4584 &  n_33069;
assign n_33071 = ~n_4578 &  n_33070;
assign n_33072 = ~n_4572 &  n_33071;
assign n_33073 = ~n_4566 &  n_33072;
assign n_33074 = ~n_4560 &  n_33073;
assign n_33075 = ~n_4554 &  n_33074;
assign n_33076 = ~n_4548 &  n_33075;
assign n_33077 = ~n_4542 &  n_33076;
assign n_33078 = ~n_4536 &  n_33077;
assign n_33079 = ~n_4530 &  n_33078;
assign n_33080 = ~n_4524 &  n_33079;
assign n_33081 = ~n_4518 &  n_33080;
assign n_33082 = ~n_4512 &  n_33081;
assign n_33083 = ~n_4506 &  n_33082;
assign n_33084 = ~n_4500 &  n_33083;
assign n_33085 = ~n_4494 &  n_33084;
assign n_33086 = ~n_4488 &  n_33085;
assign n_33087 = ~n_4482 &  n_33086;
assign n_33088 = ~n_4476 &  n_33087;
assign n_33089 = ~n_4470 &  n_33088;
assign n_33090 = ~n_4464 &  n_33089;
assign n_33091 = ~n_4458 &  n_33090;
assign n_33092 = ~n_4452 &  n_33091;
assign n_33093 = ~n_4444 &  n_33092;
assign n_33094 = ~n_4438 &  n_33093;
assign n_33095 = ~n_4432 &  n_33094;
assign n_33096 = ~n_4426 &  n_33095;
assign n_33097 = ~n_4420 &  n_33096;
assign n_33098 = ~n_4414 &  n_33097;
assign n_33099 = ~n_4408 &  n_33098;
assign n_33100 = ~n_4402 &  n_33099;
assign n_33101 = ~n_4396 &  n_33100;
assign n_33102 = ~n_4390 &  n_33101;
assign n_33103 = ~n_4384 &  n_33102;
assign n_33104 = ~n_4378 &  n_33103;
assign n_33105 = ~n_4372 &  n_33104;
assign n_33106 = ~n_4366 &  n_33105;
assign n_33107 = ~n_4360 &  n_33106;
assign n_33108 = ~n_4354 &  n_33107;
assign n_33109 = ~n_4348 &  n_33108;
assign n_33110 = ~n_4342 &  n_33109;
assign n_33111 = ~n_4336 &  n_33110;
assign n_33112 = ~n_4330 &  n_33111;
assign n_33113 = ~n_4324 &  n_33112;
assign n_33114 = ~n_4318 &  n_33113;
assign n_33115 = ~n_4312 &  n_33114;
assign n_33116 = ~n_4306 &  n_33115;
assign n_33117 = ~n_4300 &  n_33116;
assign n_33118 = ~n_4294 &  n_33117;
assign n_33119 = ~n_4288 &  n_33118;
assign n_33120 = ~n_4282 &  n_33119;
assign n_33121 = ~n_4276 &  n_33120;
assign n_33122 = ~n_4270 &  n_33121;
assign n_33123 = ~n_4264 &  n_33122;
assign n_33124 = ~n_4258 &  n_33123;
assign n_33125 = ~n_4250 &  n_33124;
assign n_33126 = ~n_4244 &  n_33125;
assign n_33127 = ~n_4238 &  n_33126;
assign n_33128 = ~n_4232 &  n_33127;
assign n_33129 = ~n_4226 &  n_33128;
assign n_33130 = ~n_4220 &  n_33129;
assign n_33131 = ~n_4214 &  n_33130;
assign n_33132 = ~n_4208 &  n_33131;
assign n_33133 = ~n_4202 &  n_33132;
assign n_33134 = ~n_4196 &  n_33133;
assign n_33135 = ~n_4190 &  n_33134;
assign n_33136 = ~n_4184 &  n_33135;
assign n_33137 = ~n_4178 &  n_33136;
assign n_33138 = ~n_4172 &  n_33137;
assign n_33139 = ~n_4166 &  n_33138;
assign n_33140 = ~n_4160 &  n_33139;
assign n_33141 = ~n_4154 &  n_33140;
assign n_33142 = ~n_4148 &  n_33141;
assign n_33143 = ~n_4142 &  n_33142;
assign n_33144 = ~n_4136 &  n_33143;
assign n_33145 = ~n_4130 &  n_33144;
assign n_33146 = ~n_4124 &  n_33145;
assign n_33147 = ~n_4118 &  n_33146;
assign n_33148 = ~n_4112 &  n_33147;
assign n_33149 = ~n_4106 &  n_33148;
assign n_33150 = ~n_4100 &  n_33149;
assign n_33151 = ~n_4094 &  n_33150;
assign n_33152 = ~n_4088 &  n_33151;
assign n_33153 = ~n_4082 &  n_33152;
assign n_33154 = ~n_4076 &  n_33153;
assign n_33155 = ~n_4070 &  n_33154;
assign n_33156 = ~n_4064 &  n_33155;
assign n_33157 = ~n_4055 &  n_33156;
assign n_33158 = ~n_4049 &  n_33157;
assign n_33159 = ~n_4043 &  n_33158;
assign n_33160 = ~n_4037 &  n_33159;
assign n_33161 = ~n_4031 &  n_33160;
assign n_33162 = ~n_4025 &  n_33161;
assign n_33163 = ~n_4019 &  n_33162;
assign n_33164 = ~n_4013 &  n_33163;
assign n_33165 = ~n_4007 &  n_33164;
assign n_33166 = ~n_4001 &  n_33165;
assign n_33167 = ~n_3995 &  n_33166;
assign n_33168 = ~n_3989 &  n_33167;
assign n_33169 = ~n_3983 &  n_33168;
assign n_33170 = ~n_3977 &  n_33169;
assign n_33171 = ~n_3971 &  n_33170;
assign n_33172 = ~n_3965 &  n_33171;
assign n_33173 = ~n_3959 &  n_33172;
assign n_33174 = ~n_3953 &  n_33173;
assign n_33175 = ~n_3947 &  n_33174;
assign n_33176 = ~n_3941 &  n_33175;
assign n_33177 = ~n_3935 &  n_33176;
assign n_33178 = ~n_3929 &  n_33177;
assign n_33179 = ~n_3923 &  n_33178;
assign n_33180 = ~n_3917 &  n_33179;
assign n_33181 = ~n_3911 &  n_33180;
assign n_33182 = ~n_3905 &  n_33181;
assign n_33183 = ~n_3899 &  n_33182;
assign n_33184 = ~n_3893 &  n_33183;
assign n_33185 = ~n_3887 &  n_33184;
assign n_33186 = ~n_3881 &  n_33185;
assign n_33187 = ~n_3875 &  n_33186;
assign n_33188 = ~n_3869 &  n_33187;
assign n_33189 = ~n_3857 &  n_33188;
assign n_33190 = ~n_3851 &  n_33189;
assign n_33191 = ~n_3845 &  n_33190;
assign n_33192 = ~n_3839 &  n_33191;
assign n_33193 = ~n_3833 &  n_33192;
assign n_33194 = ~n_3827 &  n_33193;
assign n_33195 = ~n_3821 &  n_33194;
assign n_33196 = ~n_3815 &  n_33195;
assign n_33197 = ~n_3809 &  n_33196;
assign n_33198 = ~n_3803 &  n_33197;
assign n_33199 = ~n_3797 &  n_33198;
assign n_33200 = ~n_3791 &  n_33199;
assign n_33201 = ~n_3785 &  n_33200;
assign n_33202 = ~n_3779 &  n_33201;
assign n_33203 = ~n_3773 &  n_33202;
assign n_33204 = ~n_3767 &  n_33203;
assign n_33205 = ~n_3761 &  n_33204;
assign n_33206 = ~n_3755 &  n_33205;
assign n_33207 = ~n_3749 &  n_33206;
assign n_33208 = ~n_3743 &  n_33207;
assign n_33209 = ~n_3737 &  n_33208;
assign n_33210 = ~n_3731 &  n_33209;
assign n_33211 = ~n_3725 &  n_33210;
assign n_33212 = ~n_3719 &  n_33211;
assign n_33213 = ~n_3713 &  n_33212;
assign n_33214 = ~n_3707 &  n_33213;
assign n_33215 = ~n_3701 &  n_33214;
assign n_33216 = ~n_3695 &  n_33215;
assign n_33217 = ~n_3689 &  n_33216;
assign n_33218 = ~n_3683 &  n_33217;
assign n_33219 = ~n_3677 &  n_33218;
assign n_33220 = ~n_3671 &  n_33219;
assign n_33221 = ~n_3662 &  n_33220;
assign n_33222 = ~n_3656 &  n_33221;
assign n_33223 = ~n_3650 &  n_33222;
assign n_33224 = ~n_3644 &  n_33223;
assign n_33225 = ~n_3638 &  n_33224;
assign n_33226 = ~n_3632 &  n_33225;
assign n_33227 = ~n_3626 &  n_33226;
assign n_33228 = ~n_3620 &  n_33227;
assign n_33229 = ~n_3614 &  n_33228;
assign n_33230 = ~n_3608 &  n_33229;
assign n_33231 = ~n_3602 &  n_33230;
assign n_33232 = ~n_3596 &  n_33231;
assign n_33233 = ~n_3590 &  n_33232;
assign n_33234 = ~n_3584 &  n_33233;
assign n_33235 = ~n_3578 &  n_33234;
assign n_33236 = ~n_3572 &  n_33235;
assign n_33237 = ~n_3566 &  n_33236;
assign n_33238 = ~n_3560 &  n_33237;
assign n_33239 = ~n_3554 &  n_33238;
assign n_33240 = ~n_3548 &  n_33239;
assign n_33241 = ~n_3542 &  n_33240;
assign n_33242 = ~n_3536 &  n_33241;
assign n_33243 = ~n_3530 &  n_33242;
assign n_33244 = ~n_3524 &  n_33243;
assign n_33245 = ~n_3518 &  n_33244;
assign n_33246 = ~n_3512 &  n_33245;
assign n_33247 = ~n_3506 &  n_33246;
assign n_33248 = ~n_3500 &  n_33247;
assign n_33249 = ~n_3494 &  n_33248;
assign n_33250 = ~n_3488 &  n_33249;
assign n_33251 = ~n_3482 &  n_33250;
assign n_33252 = ~n_3476 &  n_33251;
assign n_33253 = ~n_3468 &  n_33252;
assign n_33254 = ~n_3462 &  n_33253;
assign n_33255 = ~n_3456 &  n_33254;
assign n_33256 = ~n_3450 &  n_33255;
assign n_33257 = ~n_3444 &  n_33256;
assign n_33258 = ~n_3438 &  n_33257;
assign n_33259 = ~n_3432 &  n_33258;
assign n_33260 = ~n_3426 &  n_33259;
assign n_33261 = ~n_3420 &  n_33260;
assign n_33262 = ~n_3414 &  n_33261;
assign n_33263 = ~n_3408 &  n_33262;
assign n_33264 = ~n_3402 &  n_33263;
assign n_33265 = ~n_3396 &  n_33264;
assign n_33266 = ~n_3390 &  n_33265;
assign n_33267 = ~n_3384 &  n_33266;
assign n_33268 = ~n_3378 &  n_33267;
assign n_33269 = ~n_3372 &  n_33268;
assign n_33270 = ~n_3366 &  n_33269;
assign n_33271 = ~n_3360 &  n_33270;
assign n_33272 = ~n_3354 &  n_33271;
assign n_33273 = ~n_3348 &  n_33272;
assign n_33274 = ~n_3342 &  n_33273;
assign n_33275 = ~n_3336 &  n_33274;
assign n_33276 = ~n_3330 &  n_33275;
assign n_33277 = ~n_3324 &  n_33276;
assign n_33278 = ~n_3318 &  n_33277;
assign n_33279 = ~n_3312 &  n_33278;
assign n_33280 = ~n_3306 &  n_33279;
assign n_33281 = ~n_3300 &  n_33280;
assign n_33282 = ~n_3294 &  n_33281;
assign n_33283 = ~n_3288 &  n_33282;
assign n_33284 = ~n_3282 &  n_33283;
assign n_33285 = ~n_3274 &  n_33284;
assign n_33286 = ~n_3268 &  n_33285;
assign n_33287 = ~n_3262 &  n_33286;
assign n_33288 = ~n_3256 &  n_33287;
assign n_33289 = ~n_3250 &  n_33288;
assign n_33290 = ~n_3244 &  n_33289;
assign n_33291 = ~n_3238 &  n_33290;
assign n_33292 = ~n_3232 &  n_33291;
assign n_33293 = ~n_3226 &  n_33292;
assign n_33294 = ~n_3220 &  n_33293;
assign n_33295 = ~n_3214 &  n_33294;
assign n_33296 = ~n_3208 &  n_33295;
assign n_33297 = ~n_3202 &  n_33296;
assign n_33298 = ~n_3196 &  n_33297;
assign n_33299 = ~n_3190 &  n_33298;
assign n_33300 = ~n_3184 &  n_33299;
assign n_33301 = ~n_3178 &  n_33300;
assign n_33302 = ~n_3172 &  n_33301;
assign n_33303 = ~n_3166 &  n_33302;
assign n_33304 = ~n_3160 &  n_33303;
assign n_33305 = ~n_3154 &  n_33304;
assign n_33306 = ~n_3148 &  n_33305;
assign n_33307 = ~n_3142 &  n_33306;
assign n_33308 = ~n_3136 &  n_33307;
assign n_33309 = ~n_3130 &  n_33308;
assign n_33310 = ~n_3124 &  n_33309;
assign n_33311 = ~n_3118 &  n_33310;
assign n_33312 = ~n_3112 &  n_33311;
assign n_33313 = ~n_3106 &  n_33312;
assign n_33314 = ~n_3100 &  n_33313;
assign n_33315 = ~n_3094 &  n_33314;
assign n_33316 = ~n_3088 &  n_33315;
assign n_33317 = ~n_3080 &  n_33316;
assign n_33318 = ~n_3074 &  n_33317;
assign n_33319 = ~n_3068 &  n_33318;
assign n_33320 = ~n_3062 &  n_33319;
assign n_33321 = ~n_3056 &  n_33320;
assign n_33322 = ~n_3050 &  n_33321;
assign n_33323 = ~n_3044 &  n_33322;
assign n_33324 = ~n_3038 &  n_33323;
assign n_33325 = ~n_3032 &  n_33324;
assign n_33326 = ~n_3026 &  n_33325;
assign n_33327 = ~n_3020 &  n_33326;
assign n_33328 = ~n_3014 &  n_33327;
assign n_33329 = ~n_3008 &  n_33328;
assign n_33330 = ~n_3002 &  n_33329;
assign n_33331 = ~n_2996 &  n_33330;
assign n_33332 = ~n_2990 &  n_33331;
assign n_33333 = ~n_2984 &  n_33332;
assign n_33334 = ~n_2978 &  n_33333;
assign n_33335 = ~n_2972 &  n_33334;
assign n_33336 = ~n_2966 &  n_33335;
assign n_33337 = ~n_2960 &  n_33336;
assign n_33338 = ~n_2954 &  n_33337;
assign n_33339 = ~n_2948 &  n_33338;
assign n_33340 = ~n_2942 &  n_33339;
assign n_33341 = ~n_2936 &  n_33340;
assign n_33342 = ~n_2930 &  n_33341;
assign n_33343 = ~n_2924 &  n_33342;
assign n_33344 = ~n_2918 &  n_33343;
assign n_33345 = ~n_2912 &  n_33344;
assign n_33346 = ~n_2906 &  n_33345;
assign n_33347 = ~n_2900 &  n_33346;
assign n_33348 = ~n_2894 &  n_33347;
assign n_33349 = ~n_2885 &  n_33348;
assign n_33350 = ~n_2879 &  n_33349;
assign n_33351 = ~n_2873 &  n_33350;
assign n_33352 = ~n_2867 &  n_33351;
assign n_33353 = ~n_2861 &  n_33352;
assign n_33354 = ~n_2855 &  n_33353;
assign n_33355 = ~n_2849 &  n_33354;
assign n_33356 = ~n_2843 &  n_33355;
assign n_33357 = ~n_2837 &  n_33356;
assign n_33358 = ~n_2831 &  n_33357;
assign n_33359 = ~n_2825 &  n_33358;
assign n_33360 = ~n_2819 &  n_33359;
assign n_33361 = ~n_2813 &  n_33360;
assign n_33362 = ~n_2807 &  n_33361;
assign n_33363 = ~n_2801 &  n_33362;
assign n_33364 = ~n_2795 &  n_33363;
assign n_33365 = ~n_2789 &  n_33364;
assign n_33366 = ~n_2783 &  n_33365;
assign n_33367 = ~n_2777 &  n_33366;
assign n_33368 = ~n_2771 &  n_33367;
assign n_33369 = ~n_2765 &  n_33368;
assign n_33370 = ~n_2759 &  n_33369;
assign n_33371 = ~n_2753 &  n_33370;
assign n_33372 = ~n_2747 &  n_33371;
assign n_33373 = ~n_2741 &  n_33372;
assign n_33374 = ~n_2735 &  n_33373;
assign n_33375 = ~n_2729 &  n_33374;
assign n_33376 = ~n_2723 &  n_33375;
assign n_33377 = ~n_2717 &  n_33376;
assign n_33378 = ~n_2711 &  n_33377;
assign n_33379 = ~n_2705 &  n_33378;
assign n_33380 = ~n_2699 &  n_33379;
assign n_33381 = ~n_2692 &  n_33380;
assign n_33382 = ~n_2686 &  n_33381;
assign n_33383 = ~n_2680 &  n_33382;
assign n_33384 = ~n_2674 &  n_33383;
assign n_33385 = ~n_2668 &  n_33384;
assign n_33386 = ~n_2662 &  n_33385;
assign n_33387 = ~n_2656 &  n_33386;
assign n_33388 = ~n_2650 &  n_33387;
assign n_33389 = ~n_2644 &  n_33388;
assign n_33390 = ~n_2638 &  n_33389;
assign n_33391 = ~n_2632 &  n_33390;
assign n_33392 = ~n_2626 &  n_33391;
assign n_33393 = ~n_2620 &  n_33392;
assign n_33394 = ~n_2614 &  n_33393;
assign n_33395 = ~n_2608 &  n_33394;
assign n_33396 = ~n_2602 &  n_33395;
assign n_33397 = ~n_2596 &  n_33396;
assign n_33398 = ~n_2590 &  n_33397;
assign n_33399 = ~n_2584 &  n_33398;
assign n_33400 = ~n_2578 &  n_33399;
assign n_33401 = ~n_2572 &  n_33400;
assign n_33402 = ~n_2566 &  n_33401;
assign n_33403 = ~n_2560 &  n_33402;
assign n_33404 = ~n_2554 &  n_33403;
assign n_33405 = ~n_2548 &  n_33404;
assign n_33406 = ~n_2542 &  n_33405;
assign n_33407 = ~n_2536 &  n_33406;
assign n_33408 = ~n_2530 &  n_33407;
assign n_33409 = ~n_2524 &  n_33408;
assign n_33410 = ~n_2518 &  n_33409;
assign n_33411 = ~n_2512 &  n_33410;
assign n_33412 = ~n_2506 &  n_33411;
assign n_33413 = ~n_2498 &  n_33412;
assign n_33414 = ~n_2492 &  n_33413;
assign n_33415 = ~n_2486 &  n_33414;
assign n_33416 = ~n_2480 &  n_33415;
assign n_33417 = ~n_2474 &  n_33416;
assign n_33418 = ~n_2468 &  n_33417;
assign n_33419 = ~n_2462 &  n_33418;
assign n_33420 = ~n_2456 &  n_33419;
assign n_33421 = ~n_2450 &  n_33420;
assign n_33422 = ~n_2444 &  n_33421;
assign n_33423 = ~n_2438 &  n_33422;
assign n_33424 = ~n_2432 &  n_33423;
assign n_33425 = ~n_2426 &  n_33424;
assign n_33426 = ~n_2420 &  n_33425;
assign n_33427 = ~n_2414 &  n_33426;
assign n_33428 = ~n_2408 &  n_33427;
assign n_33429 = ~n_2402 &  n_33428;
assign n_33430 = ~n_2396 &  n_33429;
assign n_33431 = ~n_2390 &  n_33430;
assign n_33432 = ~n_2384 &  n_33431;
assign n_33433 = ~n_2378 &  n_33432;
assign n_33434 = ~n_2372 &  n_33433;
assign n_33435 = ~n_2366 &  n_33434;
assign n_33436 = ~n_2360 &  n_33435;
assign n_33437 = ~n_2354 &  n_33436;
assign n_33438 = ~n_2348 &  n_33437;
assign n_33439 = ~n_2342 &  n_33438;
assign n_33440 = ~n_2336 &  n_33439;
assign n_33441 = ~n_2330 &  n_33440;
assign n_33442 = ~n_2324 &  n_33441;
assign n_33443 = ~n_2318 &  n_33442;
assign n_33444 = ~n_2312 &  n_33443;
assign n_33445 = ~n_2294 &  n_33444;
assign n_33446 = ~n_2288 &  n_33445;
assign n_33447 = ~n_2282 &  n_33446;
assign n_33448 = ~n_2276 &  n_33447;
assign n_33449 = ~n_2270 &  n_33448;
assign n_33450 = ~n_2264 &  n_33449;
assign n_33451 = ~n_2258 &  n_33450;
assign n_33452 = ~n_2252 &  n_33451;
assign n_33453 = ~n_2246 &  n_33452;
assign n_33454 = ~n_2240 &  n_33453;
assign n_33455 = ~n_2234 &  n_33454;
assign n_33456 = ~n_2228 &  n_33455;
assign n_33457 = ~n_2222 &  n_33456;
assign n_33458 = ~n_2216 &  n_33457;
assign n_33459 = ~n_2210 &  n_33458;
assign n_33460 = ~n_2204 &  n_33459;
assign n_33461 = ~n_2198 &  n_33460;
assign n_33462 = ~n_2192 &  n_33461;
assign n_33463 = ~n_2186 &  n_33462;
assign n_33464 = ~n_2180 &  n_33463;
assign n_33465 = ~n_2174 &  n_33464;
assign n_33466 = ~n_2168 &  n_33465;
assign n_33467 = ~n_2162 &  n_33466;
assign n_33468 = ~n_2156 &  n_33467;
assign n_33469 = ~n_2150 &  n_33468;
assign n_33470 = ~n_2144 &  n_33469;
assign n_33471 = ~n_2138 &  n_33470;
assign n_33472 = ~n_2132 &  n_33471;
assign n_33473 = ~n_2126 &  n_33472;
assign n_33474 = ~n_2120 &  n_33473;
assign n_33475 = ~n_2114 &  n_33474;
assign n_33476 = ~n_2108 &  n_33475;
assign n_33477 = ~n_2099 &  n_33476;
assign n_33478 = ~n_2093 &  n_33477;
assign n_33479 = ~n_2087 &  n_33478;
assign n_33480 = ~n_2081 &  n_33479;
assign n_33481 = ~n_2075 &  n_33480;
assign n_33482 = ~n_2069 &  n_33481;
assign n_33483 = ~n_2063 &  n_33482;
assign n_33484 = ~n_2057 &  n_33483;
assign n_33485 = ~n_2051 &  n_33484;
assign n_33486 = ~n_2045 &  n_33485;
assign n_33487 = ~n_2039 &  n_33486;
assign n_33488 = ~n_2033 &  n_33487;
assign n_33489 = ~n_2027 &  n_33488;
assign n_33490 = ~n_2021 &  n_33489;
assign n_33491 = ~n_2015 &  n_33490;
assign n_33492 = ~n_2009 &  n_33491;
assign n_33493 = ~n_2003 &  n_33492;
assign n_33494 = ~n_1997 &  n_33493;
assign n_33495 = ~n_1991 &  n_33494;
assign n_33496 = ~n_1985 &  n_33495;
assign n_33497 = ~n_1979 &  n_33496;
assign n_33498 = ~n_1973 &  n_33497;
assign n_33499 = ~n_1967 &  n_33498;
assign n_33500 = ~n_1961 &  n_33499;
assign n_33501 = ~n_1955 &  n_33500;
assign n_33502 = ~n_1949 &  n_33501;
assign n_33503 = ~n_1943 &  n_33502;
assign n_33504 = ~n_1937 &  n_33503;
assign n_33505 = ~n_1931 &  n_33504;
assign n_33506 = ~n_1925 &  n_33505;
assign n_33507 = ~n_1919 &  n_33506;
assign n_33508 = ~n_1913 &  n_33507;
assign n_33509 = ~n_1902 &  n_33508;
assign n_33510 = ~n_1896 &  n_33509;
assign n_33511 = ~n_1890 &  n_33510;
assign n_33512 = ~n_1884 &  n_33511;
assign n_33513 = ~n_1878 &  n_33512;
assign n_33514 = ~n_1872 &  n_33513;
assign n_33515 = ~n_1866 &  n_33514;
assign n_33516 = ~n_1860 &  n_33515;
assign n_33517 = ~n_1854 &  n_33516;
assign n_33518 = ~n_1848 &  n_33517;
assign n_33519 = ~n_1842 &  n_33518;
assign n_33520 = ~n_1836 &  n_33519;
assign n_33521 = ~n_1830 &  n_33520;
assign n_33522 = ~n_1824 &  n_33521;
assign n_33523 = ~n_1818 &  n_33522;
assign n_33524 = ~n_1812 &  n_33523;
assign n_33525 = ~n_1806 &  n_33524;
assign n_33526 = ~n_1800 &  n_33525;
assign n_33527 = ~n_1794 &  n_33526;
assign n_33528 = ~n_1788 &  n_33527;
assign n_33529 = ~n_1782 &  n_33528;
assign n_33530 = ~n_1776 &  n_33529;
assign n_33531 = ~n_1770 &  n_33530;
assign n_33532 = ~n_1764 &  n_33531;
assign n_33533 = ~n_1758 &  n_33532;
assign n_33534 = ~n_1752 &  n_33533;
assign n_33535 = ~n_1746 &  n_33534;
assign n_33536 = ~n_1740 &  n_33535;
assign n_33537 = ~n_1734 &  n_33536;
assign n_33538 = ~n_1728 &  n_33537;
assign n_33539 = ~n_1722 &  n_33538;
assign n_33540 = ~n_1716 &  n_33539;
assign n_33541 = ~n_1705 &  n_33540;
assign n_33542 = ~n_1699 &  n_33541;
assign n_33543 = ~n_1693 &  n_33542;
assign n_33544 = ~n_1687 &  n_33543;
assign n_33545 = ~n_1681 &  n_33544;
assign n_33546 = ~n_1675 &  n_33545;
assign n_33547 = ~n_1669 &  n_33546;
assign n_33548 = ~n_1663 &  n_33547;
assign n_33549 = ~n_1657 &  n_33548;
assign n_33550 = ~n_1651 &  n_33549;
assign n_33551 = ~n_1645 &  n_33550;
assign n_33552 = ~n_1639 &  n_33551;
assign n_33553 = ~n_1633 &  n_33552;
assign n_33554 = ~n_1627 &  n_33553;
assign n_33555 = ~n_1621 &  n_33554;
assign n_33556 = ~n_1615 &  n_33555;
assign n_33557 = ~n_1609 &  n_33556;
assign n_33558 = ~n_1603 &  n_33557;
assign n_33559 = ~n_1597 &  n_33558;
assign n_33560 = ~n_1591 &  n_33559;
assign n_33561 = ~n_1585 &  n_33560;
assign n_33562 = ~n_1579 &  n_33561;
assign n_33563 = ~n_1573 &  n_33562;
assign n_33564 = ~n_1567 &  n_33563;
assign n_33565 = ~n_1561 &  n_33564;
assign n_33566 = ~n_1555 &  n_33565;
assign n_33567 = ~n_1549 &  n_33566;
assign n_33568 = ~n_1543 &  n_33567;
assign n_33569 = ~n_1537 &  n_33568;
assign n_33570 = ~n_1531 &  n_33569;
assign n_33571 = ~n_1525 &  n_33570;
assign n_33572 = ~n_1519 &  n_33571;
assign n_33573 = ~n_1509 &  n_33572;
assign n_33574 = ~n_1503 &  n_33573;
assign n_33575 = ~n_1497 &  n_33574;
assign n_33576 = ~n_1491 &  n_33575;
assign n_33577 = ~n_1485 &  n_33576;
assign n_33578 = ~n_1479 &  n_33577;
assign n_33579 = ~n_1473 &  n_33578;
assign n_33580 = ~n_1467 &  n_33579;
assign n_33581 = ~n_1461 &  n_33580;
assign n_33582 = ~n_1455 &  n_33581;
assign n_33583 = ~n_1449 &  n_33582;
assign n_33584 = ~n_1443 &  n_33583;
assign n_33585 = ~n_1437 &  n_33584;
assign n_33586 = ~n_1431 &  n_33585;
assign n_33587 = ~n_1425 &  n_33586;
assign n_33588 = ~n_1419 &  n_33587;
assign n_33589 = ~n_1413 &  n_33588;
assign n_33590 = ~n_1407 &  n_33589;
assign n_33591 = ~n_1401 &  n_33590;
assign n_33592 = ~n_1395 &  n_33591;
assign n_33593 = ~n_1389 &  n_33592;
assign n_33594 = ~n_1383 &  n_33593;
assign n_33595 = ~n_1377 &  n_33594;
assign n_33596 = ~n_1371 &  n_33595;
assign n_33597 = ~n_1365 &  n_33596;
assign n_33598 = ~n_1359 &  n_33597;
assign n_33599 = ~n_1353 &  n_33598;
assign n_33600 = ~n_1347 &  n_33599;
assign n_33601 = ~n_1341 &  n_33600;
assign n_33602 = ~n_1335 &  n_33601;
assign n_33603 = ~n_1329 &  n_33602;
assign n_33604 = ~n_1323 &  n_33603;
assign n_33605 = ~n_1310 &  n_33604;
assign n_33606 = ~n_1306 &  n_33605;
assign n_33607 = ~n_1302 &  n_33606;
assign n_33608 = ~n_1298 &  n_33607;
assign n_33609 = ~n_1294 &  n_33608;
assign n_33610 = ~n_1290 &  n_33609;
assign n_33611 = ~n_1286 &  n_33610;
assign n_33612 = ~n_1282 &  n_33611;
assign n_33613 = ~n_1278 &  n_33612;
assign n_33614 = ~n_1274 &  n_33613;
assign n_33615 = ~n_1270 &  n_33614;
assign n_33616 = ~n_1266 &  n_33615;
assign n_33617 = ~n_1262 &  n_33616;
assign n_33618 = ~n_1258 &  n_33617;
assign n_33619 = ~n_1254 &  n_33618;
assign n_33620 = ~n_1250 &  n_33619;
assign n_33621 = ~n_1246 &  n_33620;
assign n_33622 = ~n_1242 &  n_33621;
assign n_33623 = ~n_1238 &  n_33622;
assign n_33624 = ~n_1234 &  n_33623;
assign n_33625 = ~n_1230 &  n_33624;
assign n_33626 = ~n_1226 &  n_33625;
assign n_33627 = ~n_1222 &  n_33626;
assign n_33628 = ~n_1218 &  n_33627;
assign n_33629 = ~n_1214 &  n_33628;
assign n_33630 = ~n_1210 &  n_33629;
assign n_33631 = ~n_1206 &  n_33630;
assign n_33632 = ~n_1202 &  n_33631;
assign n_33633 = ~n_1198 &  n_33632;
assign n_33634 = ~n_1194 &  n_33633;
assign n_33635 = ~n_1190 &  n_33634;
assign n_33636 = ~n_1186 &  n_33635;
assign n_33637 = ~n_1176 &  n_33636;
assign n_33638 = ~n_1170 &  n_33637;
assign n_33639 = ~n_1164 &  n_33638;
assign n_33640 = ~n_1158 &  n_33639;
assign n_33641 = ~n_1152 &  n_33640;
assign n_33642 = ~n_1146 &  n_33641;
assign n_33643 = ~n_1140 &  n_33642;
assign n_33644 = ~n_1134 &  n_33643;
assign n_33645 = ~n_1128 &  n_33644;
assign n_33646 = ~n_1122 &  n_33645;
assign n_33647 = ~n_1116 &  n_33646;
assign n_33648 = ~n_1110 &  n_33647;
assign n_33649 = ~n_1104 &  n_33648;
assign n_33650 = ~n_1098 &  n_33649;
assign n_33651 = ~n_1092 &  n_33650;
assign n_33652 = ~n_1086 &  n_33651;
assign n_33653 = ~n_1080 &  n_33652;
assign n_33654 = ~n_1074 &  n_33653;
assign n_33655 = ~n_1068 &  n_33654;
assign n_33656 = ~n_1062 &  n_33655;
assign n_33657 = ~n_1056 &  n_33656;
assign n_33658 = ~n_1050 &  n_33657;
assign n_33659 = ~n_1044 &  n_33658;
assign n_33660 = ~n_1038 &  n_33659;
assign n_33661 = ~n_1032 &  n_33660;
assign n_33662 = ~n_1026 &  n_33661;
assign n_33663 = ~n_1020 &  n_33662;
assign n_33664 = ~n_1014 &  n_33663;
assign n_33665 = ~n_1008 &  n_33664;
assign n_33666 = ~n_1002 &  n_33665;
assign n_33667 = ~n_996 &  n_33666;
assign n_33668 = ~n_990 &  n_33667;
assign n_33669 = ~n_978 &  n_33668;
assign n_33670 = ~n_972 &  n_33669;
assign n_33671 = ~n_966 &  n_33670;
assign n_33672 = ~n_960 &  n_33671;
assign n_33673 = ~n_954 &  n_33672;
assign n_33674 = ~n_948 &  n_33673;
assign n_33675 = ~n_942 &  n_33674;
assign n_33676 = ~n_936 &  n_33675;
assign n_33677 = ~n_930 &  n_33676;
assign n_33678 = ~n_924 &  n_33677;
assign n_33679 = ~n_918 &  n_33678;
assign n_33680 = ~n_912 &  n_33679;
assign n_33681 = ~n_906 &  n_33680;
assign n_33682 = ~n_900 &  n_33681;
assign n_33683 = ~n_894 &  n_33682;
assign n_33684 = ~n_888 &  n_33683;
assign n_33685 = ~n_882 &  n_33684;
assign n_33686 = ~n_876 &  n_33685;
assign n_33687 = ~n_870 &  n_33686;
assign n_33688 = ~n_864 &  n_33687;
assign n_33689 = ~n_858 &  n_33688;
assign n_33690 = ~n_852 &  n_33689;
assign n_33691 = ~n_846 &  n_33690;
assign n_33692 = ~n_840 &  n_33691;
assign n_33693 = ~n_834 &  n_33692;
assign n_33694 = ~n_828 &  n_33693;
assign n_33695 = ~n_822 &  n_33694;
assign n_33696 = ~n_816 &  n_33695;
assign n_33697 = ~n_810 &  n_33696;
assign n_33698 = ~n_804 &  n_33697;
assign n_33699 = ~n_798 &  n_33698;
assign n_33700 = ~n_792 &  n_33699;
assign n_33701 = ~n_781 &  n_33700;
assign n_33702 = ~n_775 &  n_33701;
assign n_33703 = ~n_769 &  n_33702;
assign n_33704 = ~n_763 &  n_33703;
assign n_33705 = ~n_757 &  n_33704;
assign n_33706 = ~n_751 &  n_33705;
assign n_33707 = ~n_745 &  n_33706;
assign n_33708 = ~n_739 &  n_33707;
assign n_33709 = ~n_733 &  n_33708;
assign n_33710 = ~n_727 &  n_33709;
assign n_33711 = ~n_721 &  n_33710;
assign n_33712 = ~n_715 &  n_33711;
assign n_33713 = ~n_709 &  n_33712;
assign n_33714 = ~n_703 &  n_33713;
assign n_33715 = ~n_697 &  n_33714;
assign n_33716 = ~n_691 &  n_33715;
assign n_33717 = ~n_685 &  n_33716;
assign n_33718 = ~n_679 &  n_33717;
assign n_33719 = ~n_673 &  n_33718;
assign n_33720 = ~n_667 &  n_33719;
assign n_33721 = ~n_661 &  n_33720;
assign n_33722 = ~n_655 &  n_33721;
assign n_33723 = ~n_649 &  n_33722;
assign n_33724 = ~n_643 &  n_33723;
assign n_33725 = ~n_637 &  n_33724;
assign n_33726 = ~n_631 &  n_33725;
assign n_33727 = ~n_625 &  n_33726;
assign n_33728 = ~n_619 &  n_33727;
assign n_33729 = ~n_613 &  n_33728;
assign n_33730 = ~n_607 &  n_33729;
assign n_33731 = ~n_601 &  n_33730;
assign n_33732 = ~n_595 &  n_33731;
assign n_33733 = ~n_584 &  n_33732;
assign n_33734 = ~n_578 &  n_33733;
assign n_33735 = ~n_572 &  n_33734;
assign n_33736 = ~n_566 &  n_33735;
assign n_33737 = ~n_560 &  n_33736;
assign n_33738 = ~n_554 &  n_33737;
assign n_33739 = ~n_548 &  n_33738;
assign n_33740 = ~n_542 &  n_33739;
assign n_33741 = ~n_536 &  n_33740;
assign n_33742 = ~n_530 &  n_33741;
assign n_33743 = ~n_524 &  n_33742;
assign n_33744 = ~n_518 &  n_33743;
assign n_33745 = ~n_512 &  n_33744;
assign n_33746 = ~n_506 &  n_33745;
assign n_33747 = ~n_500 &  n_33746;
assign n_33748 = ~n_494 &  n_33747;
assign n_33749 = ~n_488 &  n_33748;
assign n_33750 = ~n_482 &  n_33749;
assign n_33751 = ~n_476 &  n_33750;
assign n_33752 = ~n_470 &  n_33751;
assign n_33753 = ~n_464 &  n_33752;
assign n_33754 = ~n_458 &  n_33753;
assign n_33755 = ~n_452 &  n_33754;
assign n_33756 = ~n_446 &  n_33755;
assign n_33757 = ~n_440 &  n_33756;
assign n_33758 = ~n_434 &  n_33757;
assign n_33759 = ~n_428 &  n_33758;
assign n_33760 = ~n_422 &  n_33759;
assign n_33761 = ~n_416 &  n_33760;
assign n_33762 = ~n_410 &  n_33761;
assign n_33763 = ~n_404 &  n_33762;
assign n_33764 = ~n_398 &  n_33763;
assign n_33765 = ~n_384 &  n_33764;
assign n_33766 = ~n_378 &  n_33765;
assign n_33767 = ~n_372 &  n_33766;
assign n_33768 = ~n_366 &  n_33767;
assign n_33769 = ~n_360 &  n_33768;
assign n_33770 = ~n_354 &  n_33769;
assign n_33771 = ~n_348 &  n_33770;
assign n_33772 = ~n_342 &  n_33771;
assign n_33773 = ~n_336 &  n_33772;
assign n_33774 = ~n_330 &  n_33773;
assign n_33775 = ~n_324 &  n_33774;
assign n_33776 = ~n_318 &  n_33775;
assign n_33777 = ~n_312 &  n_33776;
assign n_33778 = ~n_306 &  n_33777;
assign n_33779 = ~n_300 &  n_33778;
assign n_33780 = ~n_294 &  n_33779;
assign n_33781 = ~n_288 &  n_33780;
assign n_33782 = ~n_282 &  n_33781;
assign n_33783 = ~n_276 &  n_33782;
assign n_33784 = ~n_270 &  n_33783;
assign n_33785 = ~n_264 &  n_33784;
assign n_33786 = ~n_258 &  n_33785;
assign n_33787 = ~n_252 &  n_33786;
assign n_33788 = ~n_246 &  n_33787;
assign n_33789 = ~n_240 &  n_33788;
assign n_33790 = ~n_234 &  n_33789;
assign n_33791 = ~n_228 &  n_33790;
assign n_33792 = ~n_222 &  n_33791;
assign n_33793 = ~n_216 &  n_33792;
assign n_33794 = ~n_210 &  n_33793;
assign n_33795 = ~n_204 &  n_33794;
assign n_33796 = ~n_198 &  n_33795;
assign n_33797 = ~n_183 &  n_33796;
assign n_33798 = ~n_177 &  n_33797;
assign n_33799 = ~n_171 &  n_33798;
assign n_33800 = ~n_165 &  n_33799;
assign n_33801 = ~n_159 &  n_33800;
assign n_33802 = ~n_153 &  n_33801;
assign n_33803 = ~n_147 &  n_33802;
assign n_33804 = ~n_141 &  n_33803;
assign n_33805 = ~n_135 &  n_33804;
assign n_33806 = ~n_129 &  n_33805;
assign n_33807 = ~n_123 &  n_33806;
assign n_33808 = ~n_117 &  n_33807;
assign n_33809 = ~n_111 &  n_33808;
assign n_33810 = ~n_105 &  n_33809;
assign n_33811 = ~n_99 &  n_33810;
assign n_33812 = ~n_93 &  n_33811;
assign n_33813 = ~n_87 &  n_33812;
assign n_33814 = ~n_81 &  n_33813;
assign n_33815 = ~n_75 &  n_33814;
assign n_33816 = ~n_69 &  n_33815;
assign n_33817 = ~n_63 &  n_33816;
assign n_33818 = ~n_57 &  n_33817;
assign n_33819 = ~n_51 &  n_33818;
assign n_33820 = ~n_45 &  n_33819;
assign n_33821 = ~n_39 &  n_33820;
assign n_33822 = ~n_33 &  n_33821;
assign n_33823 = ~n_27 &  n_33822;
assign n_33824 = ~n_21 &  n_33823;
assign n_33825 = ~n_15 &  n_33824;
assign o_1 = ~n_33825;
endmodule

