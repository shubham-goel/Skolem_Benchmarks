// Verilog file written by procedure Aig_ManDumpVerilog()
module test ( n0001, n0002, n0003, n0004, n0005, n0006, n0007, n0008, n0009, n0010, n0011, n0012, n0013, n0014, n0015, n0016, n0017, n0018, n0019, n0020, n0021, n0022, n0023, n0024, n0025, n0026, n0027, n0028, n0029, n0030, n0031, n0032, n0033, n0034, n0035, n0036, n0037, n0038, n0039, n0040, n0041, n0042, n0043, n0044, n0045, n0046, n0047, n0048, n0049, n0050, n0051, n0052, n0053, n0054, n0055, n0056, n0057, n0058, n0059, n0060, n0061, n0062, n0063, n0064, n0065, n0066, n0067, n0068, n0069, n0070, n0071, n0072, n0073, n0074, n0075, n0076, n0077, n0078, n0079, n0080, n0081, n0082, n0083, n0084, n0085, n0086, n0087, n0088, n0089, n0090, n0091, n0092, n0093, n0094, n0095, n0096, n0097, n0098, n0099, n0100, n0101, n0102, n0103, n0104, n0105, n0106, n0107, n0108, n0109, n0110, n0111, n0112, n0113, n0114, n0115, n0116, n0117, n0118, n0119, n0120, n0121, n0122, n0123, n0124, n0125, n0126, n0127, n0128, n0129, n0130, n0131, n0132, n0133, n0134, n0135, n0136, n0137, n0138, n0139, n0140, n0141, n0142, n0143, n0144, n0145, n0146, n0147, n0148, n0149, n0150, n0151, n0152, n0153, n0154, n0155, n0156, n0157, n0158, n0159, n0160, n0161, n0162, n0163, n0164, n0165, n0166, n0167, n0168, n0169, n0170, n0171, n0172, n0173, n0174, n0175, n0176, n0177, n0178, n0179, n0180, n0181, n0182, n0183, n0184, n0185, n0186, n0187, n0188, n0189, n0190, n0191, n0192, n0193, n0194, n0195, n0196, n0197, n0198, n0199, n0200, n0201, n0202, n0203, n0204, n0205, n0206, n0207, n0208, n0209, n0210, n0211, n0212, n0213, n0214, n0215, n0216, n0217, n0218, n0219, n0220, n0221, n0222, n0223, n0224, n0225, n0226, n0227, n0228, n0229, n0230, n0231, n0232, n0233, n0234, n0235, n0236, n0237, n0238, n0239, n0240, n0241, n0242, n0243, n0244, n0245, n0246, n0247, n0248, n0249, n0250, n0251, n0252, n0253, n0254, n0255, n0256, n0257, n0258, n0259, n0260, n0261, n0262, n0263, n0264, n0265, n0266, n0267, n0268, n0269, n0270, n0271, n0272, n0273, n0274, n0275, n0276, n0277, n0278, n0279, n0280, n0281, n0282, n0283, n0284, n0285, n0286, n0287, n0288, n0289, n0290, n0291, n0292, n0293, n0294, n0295, n0296, n0297, n0298, n0299, n0300, n0301, n0302, n0303, n0304, n0305, n0306, n0307, n0308, n0309, n0310, n0311, n0312, n0313, n0314, n0315, n0316, n0317, n0318, n0319, n0320, n0321, n0322, n0323, n0324, n0325, n0326, n0327, n0328, n0329, n0330, n0331, n0332, n0333, n0334, n0335, n0336, n0337, n0338, n0339, n0340, n0341, n0342, n0343, n0344, n0345, n0346, n0347, n0348, n0349, n0350, n0351, n0352, n0353, n0354, n0355, n0356, n0357, n0358, n0359, n0360, n0361, n0362, n0363, n0364, n0365, n0366, n0367, n0368, n0369, n0370, n0371, n0372, n0373, n0374, n0375, n0376, n0377, n0378, n0379, n0380, n0381, n0382, n0383, n0384, n0385, n0386, n0387, n0388, n0389, n0390, n0391, n0392, n0393, n0394, n0395, n0396, n0397, n0398, n0399, n0400, n0401, n0402, n0403, n0404, n0405, n0406, n0407, n0408, n0409, n0410, n0411, n0412, n0413, n0414, n0415, n0416, n0417, n0418, n0419, n0420, n0421, n0422, n0423, n0424, n0425, n0426, n0427, n0428, n0429, n0430, n0431, n0432, n0433, n0434, n0435, n0436, n0437, n0438, n0439, n0440, n0441, n0442, n0443, n0444, n0445, n0446, n0447, n0448, n0449, n0450, n0451, n0452, n0453, n0454, n0455, n0456, n0457, n0458, n0459, n0460, n0461, n0462, n0463, n0464, n0465, n0466, n0467, n0468, n0469, n0470, n0471, n0472, n0473, n0474, n0475, n0476, n0477, n0478, n0479, n0480, n0481, n0482, n0483, n0484, n0485, n0486, n0487, n0488, n0489, n0490, n0491, n0492, n0493, n0494, n0495, n0496, n0497, n0498, n0499, n0500, n0501, n0502, n0503, n0504, n0505, n0506, n0507, n0508, n0509, n0510, n0511, n0512, n0513, n0514, n0515, n0516, n0517, n0518, n0519, n0520, n0521, n0522, n0523, n0524, n0525, n0526, n0527, n0528, n0529, n0530, n0531, n0532, n0533, n0534, n0535, n0536, n0537, n0538, n0539, n0540, n0541, n0542, n0543, n0544, n0545, n0546, n0547, n0548, n0549, n0550, n0551, n0552, n0553, n0554, n0555, n0556, n0557, n0558, n0559, n0560, n0561, n0562, n0563, n0564, n0565, n0566, n0567, n0568, n0569, n0570, n0571, n0572, n0573, n0574, n0575, n0576, n0577, n0578, n0579, n0580, n0581, n0582, n0583, n0584, n0585, n0586, n0587, n0588, n0589, n0590, n0591, n0592, n0593, n0594, n0595, n0596, n0597, n0598, n0599, n0600, n0601, n0602, n0603, n0604, n0605, n0606, n0607, n0608, n0609, n0610, n0611, n0612, n0613, n0614, n0615, n0616, n0617, n0618, n0619, n0620, n0621, n0622, n0623, n0624, n0625, n0626, n0627, n0628, n0629, n0630, n0631, n0632, n0633, n0634, n0635, n0636, n0637, n0638, n0639, n0640, n0641, n0642, n0643, n0644, n0645, n0646, n0647, n0648, n0649, n0650, n0651, n0652, n0653, n0654, n0655, n0656, n0657, n0658, n0659, n0660, n0661, n0662, n0663, n0664, n0665, n0666, n0667, n0668, n0669, n0670, n0671, n0672, n0673, n0674, n0675, n0676, n0677, n0678, n0679, n0680, n0681, n0682, n0683, n0684, n0685, n0686, n0687, n0688, n0689, n0690, n0691, n0692, n0693, n0694, n0695, n0696, n0697, n0698, n0699, n0700, n0701, n0702, n0703, n0704, n0705, n0706, n0707, n0708, n0709, n0710, n0711, n0712, n0713, n0714, n0715, n0716, n0717, n0718, n0719, n0720, n0721, n0722, n0723, n0724, n0725, n0726, n0727, n0728, n0729, n0730, n0731, n0732, n0733, n0734, n0735, n0736, n0737, n0738, n0739 );
input n0001;
input n0002;
input n0003;
input n0004;
input n0005;
input n0006;
input n0007;
input n0008;
input n0009;
input n0010;
input n0011;
input n0012;
input n0013;
input n0014;
input n0015;
input n0016;
input n0017;
input n0018;
input n0019;
input n0020;
input n0021;
input n0022;
input n0023;
input n0024;
input n0025;
input n0026;
input n0027;
input n0028;
input n0029;
input n0030;
input n0031;
input n0032;
input n0033;
input n0034;
input n0035;
input n0036;
input n0037;
input n0038;
input n0039;
input n0040;
input n0041;
input n0042;
input n0043;
input n0044;
input n0045;
input n0046;
input n0047;
input n0048;
input n0049;
input n0050;
input n0051;
input n0052;
input n0053;
input n0054;
input n0055;
input n0056;
input n0057;
input n0058;
input n0059;
input n0060;
input n0061;
input n0062;
input n0063;
input n0064;
input n0065;
input n0066;
input n0067;
input n0068;
input n0069;
input n0070;
input n0071;
input n0072;
input n0073;
input n0074;
input n0075;
input n0076;
input n0077;
input n0078;
input n0079;
input n0080;
input n0081;
input n0082;
input n0083;
input n0084;
input n0085;
input n0086;
input n0087;
input n0088;
input n0089;
input n0090;
input n0091;
input n0092;
input n0093;
input n0094;
input n0095;
input n0096;
input n0097;
input n0098;
input n0099;
input n0100;
input n0101;
input n0102;
input n0103;
input n0104;
input n0105;
input n0106;
input n0107;
input n0108;
input n0109;
input n0110;
input n0111;
input n0112;
input n0113;
input n0114;
input n0115;
input n0116;
input n0117;
input n0118;
input n0119;
input n0120;
input n0121;
input n0122;
input n0123;
input n0124;
input n0125;
input n0126;
input n0127;
input n0128;
input n0129;
input n0130;
input n0131;
input n0132;
input n0133;
input n0134;
input n0135;
input n0136;
input n0137;
input n0138;
input n0139;
input n0140;
input n0141;
input n0142;
input n0143;
input n0144;
input n0145;
input n0146;
input n0147;
input n0148;
input n0149;
input n0150;
input n0151;
input n0152;
input n0153;
input n0154;
input n0155;
input n0156;
input n0157;
input n0158;
input n0159;
input n0160;
input n0161;
input n0162;
input n0163;
input n0164;
input n0165;
input n0166;
input n0167;
input n0168;
input n0169;
input n0170;
input n0171;
input n0172;
input n0173;
input n0174;
input n0175;
input n0176;
input n0177;
input n0178;
input n0179;
input n0180;
input n0181;
input n0182;
input n0183;
input n0184;
input n0185;
input n0186;
input n0187;
input n0188;
input n0189;
input n0190;
input n0191;
input n0192;
input n0193;
input n0194;
input n0195;
input n0196;
input n0197;
input n0198;
input n0199;
input n0200;
input n0201;
input n0202;
input n0203;
input n0204;
input n0205;
input n0206;
input n0207;
input n0208;
input n0209;
input n0210;
input n0211;
input n0212;
input n0213;
input n0214;
input n0215;
input n0216;
input n0217;
input n0218;
input n0219;
input n0220;
input n0221;
input n0222;
input n0223;
input n0224;
input n0225;
input n0226;
input n0227;
input n0228;
input n0229;
input n0230;
input n0231;
input n0232;
input n0233;
input n0234;
input n0235;
input n0236;
input n0237;
input n0238;
input n0239;
input n0240;
input n0241;
input n0242;
input n0243;
input n0244;
input n0245;
input n0246;
input n0247;
input n0248;
input n0249;
input n0250;
input n0251;
input n0252;
input n0253;
input n0254;
input n0255;
input n0256;
input n0257;
input n0258;
input n0259;
input n0260;
input n0261;
input n0262;
input n0263;
input n0264;
input n0265;
input n0266;
input n0267;
input n0268;
input n0269;
input n0270;
input n0271;
input n0272;
input n0273;
input n0274;
input n0275;
input n0276;
input n0277;
input n0278;
input n0279;
input n0280;
input n0281;
input n0282;
input n0283;
input n0284;
input n0285;
input n0286;
input n0287;
input n0288;
input n0289;
input n0290;
input n0291;
input n0292;
input n0293;
input n0294;
input n0295;
input n0296;
input n0297;
input n0298;
input n0299;
input n0300;
input n0301;
input n0302;
input n0303;
input n0304;
input n0305;
input n0306;
input n0307;
input n0308;
input n0309;
input n0310;
input n0311;
input n0312;
input n0313;
input n0314;
input n0315;
input n0316;
input n0317;
input n0318;
input n0319;
input n0320;
input n0321;
input n0322;
input n0323;
input n0324;
input n0325;
input n0326;
input n0327;
input n0328;
input n0329;
input n0330;
input n0331;
input n0332;
input n0333;
input n0334;
input n0335;
input n0336;
input n0337;
input n0338;
input n0339;
input n0340;
input n0341;
input n0342;
input n0343;
input n0344;
input n0345;
input n0346;
input n0347;
input n0348;
input n0349;
input n0350;
input n0351;
input n0352;
input n0353;
input n0354;
input n0355;
input n0356;
input n0357;
input n0358;
input n0359;
input n0360;
input n0361;
input n0362;
input n0363;
input n0364;
input n0365;
input n0366;
input n0367;
input n0368;
input n0369;
input n0370;
input n0371;
input n0372;
input n0373;
input n0374;
input n0375;
input n0376;
input n0377;
input n0378;
input n0379;
input n0380;
input n0381;
input n0382;
input n0383;
input n0384;
input n0385;
input n0386;
input n0387;
input n0388;
input n0389;
input n0390;
input n0391;
input n0392;
input n0393;
input n0394;
input n0395;
input n0396;
input n0397;
input n0398;
input n0399;
input n0400;
input n0401;
input n0402;
input n0403;
input n0404;
input n0405;
input n0406;
input n0407;
input n0408;
input n0409;
input n0410;
input n0411;
input n0412;
input n0413;
input n0414;
input n0415;
input n0416;
input n0417;
input n0418;
input n0419;
input n0420;
input n0421;
input n0422;
input n0423;
input n0424;
input n0425;
input n0426;
input n0427;
input n0428;
input n0429;
input n0430;
input n0431;
input n0432;
input n0433;
input n0434;
input n0435;
input n0436;
input n0437;
input n0438;
input n0439;
input n0440;
input n0441;
input n0442;
input n0443;
input n0444;
input n0445;
input n0446;
input n0447;
input n0448;
input n0449;
input n0450;
input n0451;
input n0452;
input n0453;
input n0454;
input n0455;
input n0456;
input n0457;
input n0458;
input n0459;
input n0460;
input n0461;
input n0462;
input n0463;
input n0464;
input n0465;
input n0466;
input n0467;
input n0468;
input n0469;
input n0470;
input n0471;
input n0472;
input n0473;
input n0474;
input n0475;
input n0476;
input n0477;
input n0478;
input n0479;
input n0480;
input n0481;
input n0482;
input n0483;
input n0484;
input n0485;
input n0486;
input n0487;
input n0488;
input n0489;
input n0490;
input n0491;
input n0492;
input n0493;
input n0494;
input n0495;
input n0496;
input n0497;
input n0498;
input n0499;
input n0500;
input n0501;
input n0502;
input n0503;
input n0504;
input n0505;
input n0506;
input n0507;
input n0508;
input n0509;
input n0510;
input n0511;
input n0512;
input n0513;
input n0514;
input n0515;
input n0516;
input n0517;
input n0518;
input n0519;
input n0520;
input n0521;
input n0522;
input n0523;
input n0524;
input n0525;
input n0526;
input n0527;
input n0528;
input n0529;
input n0530;
input n0531;
input n0532;
input n0533;
input n0534;
input n0535;
input n0536;
input n0537;
input n0538;
input n0539;
input n0540;
input n0541;
input n0542;
input n0543;
input n0544;
input n0545;
input n0546;
input n0547;
input n0548;
input n0549;
input n0550;
input n0551;
input n0552;
input n0553;
input n0554;
input n0555;
input n0556;
input n0557;
input n0558;
input n0559;
input n0560;
input n0561;
input n0562;
input n0563;
input n0564;
input n0565;
input n0566;
input n0567;
input n0568;
input n0569;
input n0570;
input n0571;
input n0572;
input n0573;
input n0574;
input n0575;
input n0576;
input n0577;
input n0578;
input n0579;
input n0580;
input n0581;
input n0582;
input n0583;
input n0584;
input n0585;
input n0586;
input n0587;
input n0588;
input n0589;
input n0590;
input n0591;
input n0592;
input n0593;
input n0594;
input n0595;
input n0596;
input n0597;
input n0598;
input n0599;
input n0600;
input n0601;
input n0602;
input n0603;
input n0604;
input n0605;
input n0606;
input n0607;
input n0608;
input n0609;
input n0610;
input n0611;
input n0612;
input n0613;
input n0614;
input n0615;
input n0616;
input n0617;
input n0618;
input n0619;
input n0620;
input n0621;
input n0622;
input n0623;
input n0624;
input n0625;
input n0626;
input n0627;
input n0628;
input n0629;
input n0630;
input n0631;
input n0632;
input n0633;
input n0634;
input n0635;
input n0636;
input n0637;
input n0638;
input n0639;
input n0640;
input n0641;
input n0642;
input n0643;
input n0644;
input n0645;
input n0646;
input n0647;
input n0648;
input n0649;
input n0650;
input n0651;
input n0652;
input n0653;
input n0654;
input n0655;
input n0656;
input n0657;
input n0658;
input n0659;
input n0660;
input n0661;
input n0662;
input n0663;
input n0664;
input n0665;
input n0666;
input n0667;
input n0668;
input n0669;
input n0670;
input n0671;
input n0672;
input n0673;
input n0674;
input n0675;
input n0676;
input n0677;
input n0678;
input n0679;
input n0680;
input n0681;
input n0682;
input n0683;
input n0684;
input n0685;
input n0686;
input n0687;
input n0688;
input n0689;
input n0690;
input n0691;
input n0692;
input n0693;
input n0694;
input n0695;
input n0696;
input n0697;
input n0698;
input n0699;
input n0700;
input n0701;
input n0702;
input n0703;
input n0704;
input n0705;
input n0706;
input n0707;
input n0708;
input n0709;
input n0710;
input n0711;
input n0712;
input n0713;
input n0714;
input n0715;
input n0716;
input n0717;
input n0718;
input n0719;
input n0720;
input n0721;
input n0722;
input n0723;
input n0724;
input n0725;
input n0726;
input n0727;
input n0728;
input n0729;
input n0730;
input n0731;
input n0732;
input n0733;
input n0734;
input n0735;
input n0736;
input n0737;
input n0738;
output n0739;
wire n0740;
wire n0741;
wire n0742;
wire n0743;
wire n0744;
wire n0745;
wire n0746;
wire n0747;
wire n0748;
wire n0749;
wire n0750;
wire n0751;
wire n0752;
wire n0753;
wire n0754;
wire n0755;
wire n0756;
wire n0757;
wire n0758;
wire n0759;
wire n0760;
wire n0761;
wire n0762;
wire n0763;
wire n0764;
wire n0765;
wire n0766;
wire n0767;
wire n0768;
wire n0769;
wire n0770;
wire n0771;
wire n0772;
wire n0773;
wire n0774;
wire n0775;
wire n0776;
wire n0777;
wire n0778;
wire n0779;
wire n0780;
wire n0781;
wire n0782;
wire n0783;
wire n0784;
wire n0785;
wire n0786;
wire n0787;
wire n0788;
wire n0789;
wire n0790;
wire n0791;
wire n0792;
wire n0793;
wire n0794;
wire n0795;
wire n0796;
wire n0797;
wire n0798;
wire n0799;
wire n0800;
wire n0801;
wire n0802;
wire n0803;
wire n0804;
wire n0805;
wire n0806;
wire n0807;
wire n0808;
wire n0809;
wire n0810;
wire n0811;
wire n0812;
wire n0813;
wire n0814;
wire n0815;
wire n0816;
wire n0817;
wire n0818;
wire n0819;
wire n0820;
wire n0821;
wire n0822;
wire n0823;
wire n0824;
wire n0825;
wire n0826;
wire n0827;
wire n0828;
wire n0829;
wire n0830;
wire n0831;
wire n0832;
wire n0833;
wire n0834;
wire n0835;
wire n0836;
wire n0837;
wire n0838;
wire n0839;
wire n0840;
wire n0841;
wire n0842;
wire n0843;
wire n0844;
wire n0845;
wire n0846;
wire n0847;
wire n0848;
wire n0849;
wire n0850;
wire n0851;
wire n0852;
wire n0853;
wire n0854;
wire n0855;
wire n0856;
wire n0857;
wire n0858;
wire n0859;
wire n0860;
wire n0861;
wire n0862;
wire n0863;
wire n0864;
wire n0865;
wire n0866;
wire n0867;
wire n0868;
wire n0869;
wire n0870;
wire n0871;
wire n0872;
wire n0873;
wire n0874;
wire n0875;
wire n0876;
wire n0877;
wire n0878;
wire n0879;
wire n0880;
wire n0881;
wire n0882;
wire n0883;
wire n0884;
wire n0885;
wire n0886;
wire n0887;
wire n0888;
wire n0889;
wire n0890;
wire n0891;
wire n0892;
wire n0893;
wire n0894;
wire n0895;
wire n0896;
wire n0897;
wire n0898;
wire n0899;
wire n0900;
wire n0901;
wire n0902;
wire n0903;
wire n0904;
wire n0905;
wire n0906;
wire n0907;
wire n0908;
wire n0909;
wire n0910;
wire n0911;
wire n0912;
wire n0913;
wire n0914;
wire n0915;
wire n0916;
wire n0917;
wire n0918;
wire n0919;
wire n0920;
wire n0921;
wire n0922;
wire n0923;
wire n0924;
wire n0925;
wire n0926;
wire n0927;
wire n0928;
wire n0929;
wire n0930;
wire n0931;
wire n0932;
wire n0933;
wire n0934;
wire n0935;
wire n0936;
wire n0937;
wire n0938;
wire n0939;
wire n0940;
wire n0941;
wire n0942;
wire n0943;
wire n0944;
wire n0945;
wire n0946;
wire n0947;
wire n0948;
wire n0949;
wire n0950;
wire n0951;
wire n0952;
wire n0953;
wire n0954;
wire n0955;
wire n0956;
wire n0957;
wire n0958;
wire n0959;
wire n0960;
wire n0961;
wire n0962;
wire n0963;
wire n0964;
wire n0965;
wire n0966;
wire n0967;
wire n0968;
wire n0969;
wire n0970;
wire n0971;
wire n0972;
wire n0973;
wire n0974;
wire n0975;
wire n0976;
wire n0977;
wire n0978;
wire n0979;
wire n0980;
wire n0981;
wire n0982;
wire n0983;
wire n0984;
wire n0985;
wire n0986;
wire n0987;
wire n0988;
wire n0989;
wire n0990;
wire n0991;
wire n0992;
wire n0993;
wire n0994;
wire n0995;
wire n0996;
wire n0997;
wire n0998;
wire n0999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
assign n0740 =  n0536 & ~n0738;
assign n0741 = ~n0738 & ~n0740;
assign n0742 =  n0585 & ~n0738;
assign n0743 =  n0741 & ~n0742;
assign n0744 =  n0600 & ~n0738;
assign n0745 =  n0743 & ~n0744;
assign n0746 =  n0615 & ~n0738;
assign n0747 =  n0745 & ~n0746;
assign n0748 =  n0624 & ~n0738;
assign n0749 =  n0747 & ~n0748;
assign n0750 =  n0633 & ~n0738;
assign n0751 =  n0749 & ~n0750;
assign n0752 =  n0650 & ~n0738;
assign n0753 =  n0751 & ~n0752;
assign n0754 =  n0659 & ~n0738;
assign n0755 =  n0753 & ~n0754;
assign n0756 =  n0668 & ~n0738;
assign n0757 =  n0755 & ~n0756;
assign n0758 =  n0677 & ~n0738;
assign n0759 =  n0757 & ~n0758;
assign n0760 =  n0686 & ~n0738;
assign n0761 =  n0759 & ~n0760;
assign n0762 =  n0695 & ~n0738;
assign n0763 =  n0761 & ~n0762;
assign n0764 =  n0704 & ~n0738;
assign n0765 =  n0763 & ~n0764;
assign n0766 =  n0713 & ~n0738;
assign n0767 =  n0765 & ~n0766;
assign n0768 =  n0722 & ~n0738;
assign n0769 =  n0767 & ~n0768;
assign n0770 =  n0737 & ~n0738;
assign n0771 =  n0769 & ~n0770;
assign n0772 = ~n0004 & ~n0005;
assign n0773 = ~n0006 &  n0772;
assign n0774 = ~n0003 &  n0773;
assign n0775 = ~n0002 &  n0774;
assign n0776 = ~n0001 &  n0775;
assign n0777 =  n0535 &  n0776;
assign n0778 =  n0534 &  n0777;
assign n0779 =  n0736 &  n0778;
assign n0780 = ~n0737 &  n0779;
assign n0781 =  n0771 & ~n0780;
assign n0782 =  n0729 & ~n0736;
assign n0783 =  n0781 & ~n0782;
assign n0784 =  n0735 & ~n0736;
assign n0785 =  n0783 & ~n0784;
assign n0786 =  n0526 &  n0531;
assign n0787 =  n0582 &  n0786;
assign n0788 =  n0647 &  n0787;
assign n0789 =  n0734 &  n0788;
assign n0790 = ~n0735 &  n0789;
assign n0791 =  n0785 & ~n0790;
assign n0792 =  n0733 & ~n0734;
assign n0793 =  n0791 & ~n0792;
assign n0794 =  n0336 & ~n0734;
assign n0795 =  n0793 & ~n0794;
assign n0796 =  n0337 & ~n0734;
assign n0797 =  n0795 & ~n0796;
assign n0798 =  n0338 & ~n0734;
assign n0799 =  n0797 & ~n0798;
assign n0800 =  n0339 & ~n0734;
assign n0801 =  n0799 & ~n0800;
assign n0802 =  n0731 &  n0732;
assign n0803 =  n0730 &  n0802;
assign n0804 = ~n0733 &  n0803;
assign n0805 =  n0801 & ~n0804;
assign n0806 =  n0359 & ~n0732;
assign n0807 =  n0805 & ~n0806;
assign n0808 =  n0435 & ~n0732;
assign n0809 =  n0807 & ~n0808;
assign n0810 =  n0362 & ~n0732;
assign n0811 =  n0809 & ~n0810;
assign n0812 =  n0363 & ~n0732;
assign n0813 =  n0811 & ~n0812;
assign n0814 =  n0365 & ~n0732;
assign n0815 =  n0813 & ~n0814;
assign n0816 =  n0436 & ~n0732;
assign n0817 =  n0815 & ~n0816;
assign n0818 =  n0437 & ~n0732;
assign n0819 =  n0817 & ~n0818;
assign n0820 =  n0438 & ~n0732;
assign n0821 =  n0819 & ~n0820;
assign n0822 =  n0055 & ~n0732;
assign n0823 =  n0821 & ~n0822;
assign n0824 =  n0054 & ~n0732;
assign n0825 =  n0823 & ~n0824;
assign n0826 =  n0053 & ~n0732;
assign n0827 =  n0825 & ~n0826;
assign n0828 =  n0052 & ~n0732;
assign n0829 =  n0827 & ~n0828;
assign n0830 =  n0051 & ~n0732;
assign n0831 =  n0829 & ~n0830;
assign n0832 =  n0050 & ~n0732;
assign n0833 =  n0831 & ~n0832;
assign n0834 =  n0049 & ~n0732;
assign n0835 =  n0833 & ~n0834;
assign n0836 =  n0430 & ~n0731;
assign n0837 =  n0835 & ~n0836;
assign n0838 =  n0431 & ~n0731;
assign n0839 =  n0837 & ~n0838;
assign n0840 =  n0352 & ~n0731;
assign n0841 =  n0839 & ~n0840;
assign n0842 =  n0432 & ~n0731;
assign n0843 =  n0841 & ~n0842;
assign n0844 =  n0354 & ~n0731;
assign n0845 =  n0843 & ~n0844;
assign n0846 =  n0356 & ~n0731;
assign n0847 =  n0845 & ~n0846;
assign n0848 =  n0357 & ~n0731;
assign n0849 =  n0847 & ~n0848;
assign n0850 =  n0433 & ~n0731;
assign n0851 =  n0849 & ~n0850;
assign n0852 =  n0042 & ~n0731;
assign n0853 =  n0851 & ~n0852;
assign n0854 =  n0041 & ~n0731;
assign n0855 =  n0853 & ~n0854;
assign n0856 =  n0040 & ~n0731;
assign n0857 =  n0855 & ~n0856;
assign n0858 =  n0039 & ~n0731;
assign n0859 =  n0857 & ~n0858;
assign n0860 =  n0038 & ~n0731;
assign n0861 =  n0859 & ~n0860;
assign n0862 =  n0037 & ~n0731;
assign n0863 =  n0861 & ~n0862;
assign n0864 =  n0036 & ~n0731;
assign n0865 =  n0863 & ~n0864;
assign n0866 =  n0341 & ~n0730;
assign n0867 =  n0865 & ~n0866;
assign n0868 =  n0425 & ~n0730;
assign n0869 =  n0867 & ~n0868;
assign n0870 =  n0426 & ~n0730;
assign n0871 =  n0869 & ~n0870;
assign n0872 =  n0345 & ~n0730;
assign n0873 =  n0871 & ~n0872;
assign n0874 =  n0427 & ~n0730;
assign n0875 =  n0873 & ~n0874;
assign n0876 =  n0346 & ~n0730;
assign n0877 =  n0875 & ~n0876;
assign n0878 =  n0348 & ~n0730;
assign n0879 =  n0877 & ~n0878;
assign n0880 =  n0428 & ~n0730;
assign n0881 =  n0879 & ~n0880;
assign n0882 =  n0029 & ~n0730;
assign n0883 =  n0881 & ~n0882;
assign n0884 =  n0028 & ~n0730;
assign n0885 =  n0883 & ~n0884;
assign n0886 =  n0027 & ~n0730;
assign n0887 =  n0885 & ~n0886;
assign n0888 =  n0026 & ~n0730;
assign n0889 =  n0887 & ~n0888;
assign n0890 =  n0025 & ~n0730;
assign n0891 =  n0889 & ~n0890;
assign n0892 =  n0024 & ~n0730;
assign n0893 =  n0891 & ~n0892;
assign n0894 =  n0023 & ~n0730;
assign n0895 =  n0893 & ~n0894;
assign n0896 =  n0305 &  n0306;
assign n0897 =  n0304 &  n0896;
assign n0898 =  n0303 &  n0897;
assign n0899 =  n0728 &  n0898;
assign n0900 = ~n0729 &  n0899;
assign n0901 =  n0895 & ~n0900;
assign n0902 =  n0727 & ~n0728;
assign n0903 =  n0901 & ~n0902;
assign n0904 =  n0639 & ~n0728;
assign n0905 =  n0903 & ~n0904;
assign n0906 =  n0558 & ~n0728;
assign n0907 =  n0905 & ~n0906;
assign n0908 =  n0301 & ~n0728;
assign n0909 =  n0907 & ~n0908;
assign n0910 =  n0113 &  n0114;
assign n0911 =  n0112 &  n0910;
assign n0912 =  n0111 &  n0911;
assign n0913 =  n0726 &  n0912;
assign n0914 = ~n0727 &  n0913;
assign n0915 =  n0909 & ~n0914;
assign n0916 =  n0723 & ~n0726;
assign n0917 =  n0915 & ~n0916;
assign n0918 =  n0724 & ~n0726;
assign n0919 =  n0917 & ~n0918;
assign n0920 =  n0725 & ~n0726;
assign n0921 =  n0919 & ~n0920;
assign n0922 = ~n0053 & ~n0054;
assign n0923 = ~n0055 &  n0922;
assign n0924 = ~n0052 &  n0923;
assign n0925 = ~n0050 &  n0924;
assign n0926 = ~n0051 &  n0925;
assign n0927 = ~n0049 &  n0926;
assign n0928 =  n0213 &  n0927;
assign n0929 =  n0212 &  n0928;
assign n0930 =  n0211 &  n0929;
assign n0931 =  n0140 &  n0930;
assign n0932 =  n0138 &  n0931;
assign n0933 =  n0137 &  n0932;
assign n0934 =  n0210 &  n0933;
assign n0935 =  n0134 &  n0934;
assign n0936 = ~n0725 &  n0935;
assign n0937 =  n0921 & ~n0936;
assign n0938 = ~n0038 & ~n0039;
assign n0939 = ~n0037 &  n0938;
assign n0940 = ~n0036 &  n0939;
assign n0941 = ~n0040 &  n0940;
assign n0942 = ~n0042 &  n0941;
assign n0943 = ~n0041 &  n0942;
assign n0944 =  n0208 &  n0943;
assign n0945 =  n0132 &  n0944;
assign n0946 =  n0131 &  n0945;
assign n0947 =  n0129 &  n0946;
assign n0948 =  n0207 &  n0947;
assign n0949 =  n0127 &  n0948;
assign n0950 =  n0206 &  n0949;
assign n0951 =  n0205 &  n0950;
assign n0952 = ~n0724 &  n0951;
assign n0953 =  n0937 & ~n0952;
assign n0954 = ~n0024 & ~n0025;
assign n0955 = ~n0023 &  n0954;
assign n0956 = ~n0028 &  n0955;
assign n0957 = ~n0029 &  n0956;
assign n0958 = ~n0027 &  n0957;
assign n0959 = ~n0026 &  n0958;
assign n0960 =  n0203 &  n0959;
assign n0961 =  n0123 &  n0960;
assign n0962 =  n0121 &  n0961;
assign n0963 =  n0202 &  n0962;
assign n0964 =  n0120 &  n0963;
assign n0965 =  n0201 &  n0964;
assign n0966 =  n0200 &  n0965;
assign n0967 =  n0116 &  n0966;
assign n0968 = ~n0723 &  n0967;
assign n0969 =  n0953 & ~n0968;
assign n0970 = ~n0008 &  n0772;
assign n0971 = ~n0003 &  n0970;
assign n0972 = ~n0002 &  n0971;
assign n0973 = ~n0001 &  n0972;
assign n0974 =  n0535 &  n0973;
assign n0975 =  n0534 &  n0974;
assign n0976 =  n0721 &  n0975;
assign n0977 = ~n0722 &  n0976;
assign n0978 =  n0969 & ~n0977;
assign n0979 =  n0717 & ~n0721;
assign n0980 =  n0978 & ~n0979;
assign n0981 =  n0720 & ~n0721;
assign n0982 =  n0980 & ~n0981;
assign n0983 =  n0501 &  n0531;
assign n0984 =  n0594 &  n0983;
assign n0985 =  n0500 &  n0984;
assign n0986 =  n0499 &  n0985;
assign n0987 =  n0593 &  n0986;
assign n0988 =  n0719 &  n0987;
assign n0989 =  n0718 &  n0988;
assign n0990 = ~n0720 &  n0989;
assign n0991 =  n0982 & ~n0990;
assign n0992 =  n0507 & ~n0719;
assign n0993 =  n0991 & ~n0992;
assign n0994 =  n0511 & ~n0719;
assign n0995 =  n0993 & ~n0994;
assign n0996 =  n0573 & ~n0718;
assign n0997 =  n0995 & ~n0996;
assign n0998 =  n0577 & ~n0718;
assign n0999 =  n0997 & ~n0998;
assign n1000 =  n0716 &  n0898;
assign n1001 = ~n0717 &  n1000;
assign n1002 =  n0999 & ~n1001;
assign n1003 =  n0714 & ~n0716;
assign n1004 =  n1002 & ~n1003;
assign n1005 =  n0715 & ~n0716;
assign n1006 =  n1004 & ~n1005;
assign n1007 =  n0586 & ~n0716;
assign n1008 =  n1006 & ~n1007;
assign n1009 =  n0274 & ~n0716;
assign n1010 =  n1008 & ~n1009;
assign n1011 =  n0275 & ~n0716;
assign n1012 =  n1010 & ~n1011;
assign n1013 =  n0587 & ~n0716;
assign n1014 =  n1012 & ~n1013;
assign n1015 =  n0276 & ~n0716;
assign n1016 =  n1014 & ~n1015;
assign n1017 =  n0282 &  n0286;
assign n1018 = ~n0715 &  n1017;
assign n1019 =  n1016 & ~n1018;
assign n1020 =  n0549 &  n0553;
assign n1021 = ~n0714 &  n1020;
assign n1022 =  n1019 & ~n1021;
assign n1023 = ~n0004 & ~n0007;
assign n1024 = ~n0006 &  n1023;
assign n1025 = ~n0008 &  n1024;
assign n1026 = ~n0003 &  n1025;
assign n1027 = ~n0002 &  n1026;
assign n1028 =  n0535 &  n1027;
assign n1029 =  n0534 &  n1028;
assign n1030 =  n0712 &  n1029;
assign n1031 = ~n0713 &  n1030;
assign n1032 =  n1022 & ~n1031;
assign n1033 =  n0708 & ~n0712;
assign n1034 =  n1032 & ~n1033;
assign n1035 =  n0711 & ~n0712;
assign n1036 =  n1034 & ~n1035;
assign n1037 =  n0487 &  n0531;
assign n1038 =  n0486 &  n1037;
assign n1039 =  n0485 &  n1038;
assign n1040 =  n0484 &  n1039;
assign n1041 =  n0475 &  n1040;
assign n1042 =  n0710 &  n1041;
assign n1043 =  n0709 &  n1042;
assign n1044 = ~n0711 &  n1043;
assign n1045 =  n1036 & ~n1044;
assign n1046 =  n0569 & ~n0710;
assign n1047 =  n1045 & ~n1046;
assign n1048 =  n0507 & ~n0710;
assign n1049 =  n1047 & ~n1048;
assign n1050 =  n0577 & ~n0709;
assign n1051 =  n1049 & ~n1050;
assign n1052 =  n0525 & ~n0709;
assign n1053 =  n1051 & ~n1052;
assign n1054 =  n0707 &  n0898;
assign n1055 = ~n0708 &  n1054;
assign n1056 =  n1053 & ~n1055;
assign n1057 =  n0705 & ~n0707;
assign n1058 =  n1056 & ~n1057;
assign n1059 =  n0706 & ~n0707;
assign n1060 =  n1058 & ~n1059;
assign n1061 =  n0250 & ~n0707;
assign n1062 =  n1060 & ~n1061;
assign n1063 =  n0259 & ~n0707;
assign n1064 =  n1062 & ~n1063;
assign n1065 =  n0260 & ~n0707;
assign n1066 =  n1064 & ~n1065;
assign n1067 =  n0261 & ~n0707;
assign n1068 =  n1066 & ~n1067;
assign n1069 =  n0262 & ~n0707;
assign n1070 =  n1068 & ~n1069;
assign n1071 =  n0282 &  n0545;
assign n1072 = ~n0706 &  n1071;
assign n1073 =  n1070 & ~n1072;
assign n1074 =  n0300 &  n0553;
assign n1075 = ~n0705 &  n1074;
assign n1076 =  n1073 & ~n1075;
assign n1077 = ~n0005 & ~n0007;
assign n1078 = ~n0004 &  n1077;
assign n1079 = ~n0006 &  n1078;
assign n1080 = ~n0003 &  n1079;
assign n1081 = ~n0002 &  n1080;
assign n1082 =  n0535 &  n1081;
assign n1083 =  n0534 &  n1082;
assign n1084 =  n0703 &  n1083;
assign n1085 = ~n0704 &  n1084;
assign n1086 =  n1076 & ~n1085;
assign n1087 =  n0699 & ~n0703;
assign n1088 =  n1086 & ~n1087;
assign n1089 =  n0702 & ~n0703;
assign n1090 =  n1088 & ~n1089;
assign n1091 =  n0524 &  n0531;
assign n1092 =  n0523 &  n1091;
assign n1093 =  n0518 &  n1092;
assign n1094 =  n0513 &  n1093;
assign n1095 =  n0512 &  n1094;
assign n1096 =  n0701 &  n1095;
assign n1097 =  n0700 &  n1096;
assign n1098 = ~n0702 &  n1097;
assign n1099 =  n1090 & ~n1098;
assign n1100 =  n0488 & ~n0701;
assign n1101 =  n1099 & ~n1100;
assign n1102 =  n0581 & ~n0701;
assign n1103 =  n1101 & ~n1102;
assign n1104 =  n0507 & ~n0700;
assign n1105 =  n1103 & ~n1104;
assign n1106 =  n0610 & ~n0700;
assign n1107 =  n1105 & ~n1106;
assign n1108 =  n0698 &  n0898;
assign n1109 = ~n0699 &  n1108;
assign n1110 =  n1107 & ~n1109;
assign n1111 =  n0696 & ~n0698;
assign n1112 =  n1110 & ~n1111;
assign n1113 =  n0697 & ~n0698;
assign n1114 =  n1112 & ~n1113;
assign n1115 =  n0287 & ~n0698;
assign n1116 =  n1114 & ~n1115;
assign n1117 =  n0288 & ~n0698;
assign n1118 =  n1116 & ~n1117;
assign n1119 =  n0293 & ~n0698;
assign n1120 =  n1118 & ~n1119;
assign n1121 =  n0298 & ~n0698;
assign n1122 =  n1120 & ~n1121;
assign n1123 =  n0299 & ~n0698;
assign n1124 =  n1122 & ~n1123;
assign n1125 =  n0263 &  n0557;
assign n1126 = ~n0697 &  n1125;
assign n1127 =  n1124 & ~n1126;
assign n1128 =  n0282 &  n0603;
assign n1129 = ~n0696 &  n1128;
assign n1130 =  n1127 & ~n1129;
assign n1131 = ~n0008 &  n1078;
assign n1132 = ~n0003 &  n1131;
assign n1133 = ~n0002 &  n1132;
assign n1134 =  n0535 &  n1133;
assign n1135 =  n0534 &  n1134;
assign n1136 =  n0694 &  n1135;
assign n1137 = ~n0695 &  n1136;
assign n1138 =  n1130 & ~n1137;
assign n1139 =  n0690 & ~n0694;
assign n1140 =  n1138 & ~n1139;
assign n1141 =  n0693 & ~n0694;
assign n1142 =  n1140 & ~n1141;
assign n1143 =  n0506 &  n0531;
assign n1144 =  n0505 &  n1143;
assign n1145 =  n0504 &  n1144;
assign n1146 =  n0503 &  n1145;
assign n1147 =  n0498 &  n1146;
assign n1148 =  n0692 &  n1147;
assign n1149 =  n0691 &  n1148;
assign n1150 = ~n0693 &  n1149;
assign n1151 =  n1142 & ~n1150;
assign n1152 =  n0488 & ~n0692;
assign n1153 =  n1151 & ~n1152;
assign n1154 =  n0573 & ~n0692;
assign n1155 =  n1153 & ~n1154;
assign n1156 =  n0595 & ~n0691;
assign n1157 =  n1155 & ~n1156;
assign n1158 =  n0525 & ~n0691;
assign n1159 =  n1157 & ~n1158;
assign n1160 =  n0689 &  n0898;
assign n1161 = ~n0690 &  n1160;
assign n1162 =  n1159 & ~n1161;
assign n1163 =  n0687 & ~n0689;
assign n1164 =  n1162 & ~n1163;
assign n1165 =  n0688 & ~n0689;
assign n1166 =  n1164 & ~n1165;
assign n1167 =  n0273 & ~n0689;
assign n1168 =  n1166 & ~n1167;
assign n1169 =  n0278 & ~n0689;
assign n1170 =  n1168 & ~n1169;
assign n1171 =  n0279 & ~n0689;
assign n1172 =  n1170 & ~n1171;
assign n1173 =  n0280 & ~n0689;
assign n1174 =  n1172 & ~n1173;
assign n1175 =  n0281 & ~n0689;
assign n1176 =  n1174 & ~n1175;
assign n1177 =  n0263 &  n0549;
assign n1178 = ~n0688 &  n1177;
assign n1179 =  n1176 & ~n1178;
assign n1180 =  n0300 &  n0588;
assign n1181 = ~n0687 &  n1180;
assign n1182 =  n1179 & ~n1181;
assign n1183 = ~n0004 & ~n0006;
assign n1184 = ~n0008 &  n1183;
assign n1185 = ~n0003 &  n1184;
assign n1186 = ~n0002 &  n1185;
assign n1187 = ~n0001 &  n1186;
assign n1188 =  n0535 &  n1187;
assign n1189 =  n0534 &  n1188;
assign n1190 =  n0685 &  n1189;
assign n1191 = ~n0686 &  n1190;
assign n1192 =  n1182 & ~n1191;
assign n1193 =  n0681 & ~n0685;
assign n1194 =  n1192 & ~n1193;
assign n1195 =  n0684 & ~n0685;
assign n1196 =  n1194 & ~n1195;
assign n1197 =  n0469 &  n0531;
assign n1198 =  n0576 &  n1197;
assign n1199 =  n0575 &  n1198;
assign n1200 =  n0468 &  n1199;
assign n1201 =  n0467 &  n1200;
assign n1202 =  n0683 &  n1201;
assign n1203 =  n0682 &  n1202;
assign n1204 = ~n0684 &  n1203;
assign n1205 =  n1196 & ~n1204;
assign n1206 =  n0488 & ~n0683;
assign n1207 =  n1205 & ~n1206;
assign n1208 =  n0511 & ~n0683;
assign n1209 =  n1207 & ~n1208;
assign n1210 =  n0569 & ~n0682;
assign n1211 =  n1209 & ~n1210;
assign n1212 =  n0595 & ~n0682;
assign n1213 =  n1211 & ~n1212;
assign n1214 =  n0680 &  n0898;
assign n1215 = ~n0681 &  n1214;
assign n1216 =  n1213 & ~n1215;
assign n1217 =  n0678 & ~n0680;
assign n1218 =  n1216 & ~n1217;
assign n1219 =  n0679 & ~n0680;
assign n1220 =  n1218 & ~n1219;
assign n1221 =  n0242 & ~n0680;
assign n1222 =  n1220 & ~n1221;
assign n1223 =  n0243 & ~n0680;
assign n1224 =  n1222 & ~n1223;
assign n1225 =  n0551 & ~n0680;
assign n1226 =  n1224 & ~n1225;
assign n1227 =  n0552 & ~n0680;
assign n1228 =  n1226 & ~n1227;
assign n1229 =  n0244 & ~n0680;
assign n1230 =  n1228 & ~n1229;
assign n1231 =  n0263 &  n0286;
assign n1232 = ~n0679 &  n1231;
assign n1233 =  n1230 & ~n1232;
assign n1234 =  n0545 &  n0588;
assign n1235 = ~n0678 &  n1234;
assign n1236 =  n1233 & ~n1235;
assign n1237 = ~n0005 & ~n0006;
assign n1238 = ~n0008 &  n1237;
assign n1239 = ~n0003 &  n1238;
assign n1240 = ~n0002 &  n1239;
assign n1241 = ~n0001 &  n1240;
assign n1242 =  n0535 &  n1241;
assign n1243 =  n0534 &  n1242;
assign n1244 =  n0676 &  n1243;
assign n1245 = ~n0677 &  n1244;
assign n1246 =  n1236 & ~n1245;
assign n1247 =  n0672 & ~n0676;
assign n1248 =  n1246 & ~n1247;
assign n1249 =  n0675 & ~n0676;
assign n1250 =  n1248 & ~n1249;
assign n1251 =  n0423 &  n0531;
assign n1252 =  n0510 &  n1251;
assign n1253 =  n0509 &  n1252;
assign n1254 =  n0418 &  n1253;
assign n1255 =  n0385 &  n1254;
assign n1256 =  n0674 &  n1255;
assign n1257 =  n0673 &  n1256;
assign n1258 = ~n0675 &  n1257;
assign n1259 =  n1250 & ~n1258;
assign n1260 =  n0462 & ~n0674;
assign n1261 =  n1259 & ~n1260;
assign n1262 =  n0577 & ~n0674;
assign n1263 =  n1261 & ~n1262;
assign n1264 =  n0493 & ~n0673;
assign n1265 =  n1263 & ~n1264;
assign n1266 =  n0595 & ~n0673;
assign n1267 =  n1265 & ~n1266;
assign n1268 =  n0671 &  n0898;
assign n1269 = ~n0672 &  n1268;
assign n1270 =  n1267 & ~n1269;
assign n1271 =  n0669 & ~n0671;
assign n1272 =  n1270 & ~n1271;
assign n1273 =  n0670 & ~n0671;
assign n1274 =  n1272 & ~n1273;
assign n1275 =  n0160 & ~n0671;
assign n1276 =  n1274 & ~n1275;
assign n1277 =  n0193 & ~n0671;
assign n1278 =  n1276 & ~n1277;
assign n1279 =  n0284 & ~n0671;
assign n1280 =  n1278 & ~n1279;
assign n1281 =  n0285 & ~n0671;
assign n1282 =  n1280 & ~n1281;
assign n1283 =  n0198 & ~n0671;
assign n1284 =  n1282 & ~n1283;
assign n1285 =  n0237 &  n0553;
assign n1286 = ~n0670 &  n1285;
assign n1287 =  n1284 & ~n1286;
assign n1288 =  n0268 &  n0588;
assign n1289 = ~n0669 &  n1288;
assign n1290 =  n1287 & ~n1289;
assign n1291 = ~n0006 &  n1077;
assign n1292 = ~n0008 &  n1291;
assign n1293 = ~n0002 &  n1292;
assign n1294 = ~n0001 &  n1293;
assign n1295 =  n0535 &  n1294;
assign n1296 =  n0534 &  n1295;
assign n1297 =  n0667 &  n1296;
assign n1298 = ~n0668 &  n1297;
assign n1299 =  n1290 & ~n1298;
assign n1300 =  n0663 & ~n0667;
assign n1301 =  n1299 & ~n1300;
assign n1302 =  n0666 & ~n0667;
assign n1303 =  n1301 & ~n1302;
assign n1304 =  n0452 &  n0531;
assign n1305 =  n0451 &  n1304;
assign n1306 =  n0446 &  n1305;
assign n1307 =  n0492 &  n1306;
assign n1308 =  n0490 &  n1307;
assign n1309 =  n0665 &  n1308;
assign n1310 =  n0664 &  n1309;
assign n1311 = ~n0666 &  n1310;
assign n1312 =  n1303 & ~n1311;
assign n1313 =  n0462 & ~n0665;
assign n1314 =  n1312 & ~n1313;
assign n1315 =  n0569 & ~n0665;
assign n1316 =  n1314 & ~n1315;
assign n1317 =  n0610 & ~n0664;
assign n1318 =  n1316 & ~n1317;
assign n1319 =  n0511 & ~n0664;
assign n1320 =  n1318 & ~n1319;
assign n1321 =  n0662 &  n0898;
assign n1322 = ~n0663 &  n1321;
assign n1323 =  n1320 & ~n1322;
assign n1324 =  n0660 & ~n0662;
assign n1325 =  n1323 & ~n1324;
assign n1326 =  n0661 & ~n0662;
assign n1327 =  n1325 & ~n1326;
assign n1328 =  n0265 & ~n0662;
assign n1329 =  n1327 & ~n1328;
assign n1330 =  n0267 & ~n0662;
assign n1331 =  n1329 & ~n1330;
assign n1332 =  n0221 & ~n0662;
assign n1333 =  n1331 & ~n1332;
assign n1334 =  n0226 & ~n0662;
assign n1335 =  n1333 & ~n1334;
assign n1336 =  n0227 & ~n0662;
assign n1337 =  n1335 & ~n1336;
assign n1338 =  n0237 &  n0545;
assign n1339 = ~n0661 &  n1338;
assign n1340 =  n1337 & ~n1339;
assign n1341 =  n0286 &  n0603;
assign n1342 = ~n0660 &  n1341;
assign n1343 =  n1340 & ~n1342;
assign n1344 = ~n0002 &  n1079;
assign n1345 = ~n0001 &  n1344;
assign n1346 =  n0535 &  n1345;
assign n1347 =  n0534 &  n1346;
assign n1348 =  n0658 &  n1347;
assign n1349 = ~n0659 &  n1348;
assign n1350 =  n1343 & ~n1349;
assign n1351 =  n0654 & ~n0658;
assign n1352 =  n1350 & ~n1351;
assign n1353 =  n0657 & ~n0658;
assign n1354 =  n1352 & ~n1353;
assign n1355 =  n0521 &  n0531;
assign n1356 =  n0520 &  n1355;
assign n1357 =  n0519 &  n1356;
assign n1358 =  n0609 &  n1357;
assign n1359 =  n0608 &  n1358;
assign n1360 =  n0656 &  n1359;
assign n1361 =  n0655 &  n1360;
assign n1362 = ~n0657 &  n1361;
assign n1363 =  n1354 & ~n1362;
assign n1364 =  n0493 & ~n0656;
assign n1365 =  n1363 & ~n1364;
assign n1366 =  n0525 & ~n0656;
assign n1367 =  n1365 & ~n1366;
assign n1368 =  n0569 & ~n0655;
assign n1369 =  n1367 & ~n1368;
assign n1370 =  n0581 & ~n0655;
assign n1371 =  n1369 & ~n1370;
assign n1372 =  n0653 &  n0898;
assign n1373 = ~n0654 &  n1372;
assign n1374 =  n1371 & ~n1373;
assign n1375 =  n0651 & ~n0653;
assign n1376 =  n1374 & ~n1375;
assign n1377 =  n0652 & ~n0653;
assign n1378 =  n1376 & ~n1377;
assign n1379 =  n0601 & ~n0653;
assign n1380 =  n1378 & ~n1379;
assign n1381 =  n0602 & ~n0653;
assign n1382 =  n1380 & ~n1381;
assign n1383 =  n0294 & ~n0653;
assign n1384 =  n1382 & ~n1383;
assign n1385 =  n0295 & ~n0653;
assign n1386 =  n1384 & ~n1385;
assign n1387 =  n0296 & ~n0653;
assign n1388 =  n1386 & ~n1387;
assign n1389 =  n0268 &  n0300;
assign n1390 = ~n0652 &  n1389;
assign n1391 =  n1388 & ~n1390;
assign n1392 =  n0545 &  n0557;
assign n1393 = ~n0651 &  n1392;
assign n1394 =  n1391 & ~n1393;
assign n1395 = ~n0002 &  n1131;
assign n1396 = ~n0001 &  n1395;
assign n1397 =  n0535 &  n1396;
assign n1398 =  n0534 &  n1397;
assign n1399 =  n0649 &  n1398;
assign n1400 = ~n0650 &  n1399;
assign n1401 =  n1394 & ~n1400;
assign n1402 =  n0641 & ~n0649;
assign n1403 =  n1401 & ~n1402;
assign n1404 =  n0648 & ~n0649;
assign n1405 =  n1403 & ~n1404;
assign n1406 =  n0531 &  n0647;
assign n1407 =  n0508 &  n1406;
assign n1408 =  n0574 &  n1407;
assign n1409 =  n0646 &  n1408;
assign n1410 = ~n0648 &  n1409;
assign n1411 =  n1405 & ~n1410;
assign n1412 =  n0595 & ~n0647;
assign n1413 =  n1411 & ~n1412;
assign n1414 =  n0610 & ~n0647;
assign n1415 =  n1413 & ~n1414;
assign n1416 =  n0645 & ~n0646;
assign n1417 =  n1415 & ~n1416;
assign n1418 =  n0336 & ~n0646;
assign n1419 =  n1417 & ~n1418;
assign n1420 =  n0337 & ~n0646;
assign n1421 =  n1419 & ~n1420;
assign n1422 =  n0338 & ~n0646;
assign n1423 =  n1421 & ~n1422;
assign n1424 =  n0339 & ~n0646;
assign n1425 =  n1423 & ~n1424;
assign n1426 =  n0643 &  n0644;
assign n1427 =  n0642 &  n1426;
assign n1428 = ~n0645 &  n1427;
assign n1429 =  n1425 & ~n1428;
assign n1430 =  n0396 & ~n0644;
assign n1431 =  n1429 & ~n1430;
assign n1432 =  n0412 & ~n0644;
assign n1433 =  n1431 & ~n1432;
assign n1434 =  n0397 & ~n0644;
assign n1435 =  n1433 & ~n1434;
assign n1436 =  n0413 & ~n0644;
assign n1437 =  n1435 & ~n1436;
assign n1438 =  n0414 & ~n0644;
assign n1439 =  n1437 & ~n1438;
assign n1440 =  n0398 & ~n0644;
assign n1441 =  n1439 & ~n1440;
assign n1442 =  n0415 & ~n0644;
assign n1443 =  n1441 & ~n1442;
assign n1444 =  n0399 & ~n0644;
assign n1445 =  n1443 & ~n1444;
assign n1446 =  n0073 & ~n0644;
assign n1447 =  n1445 & ~n1446;
assign n1448 =  n0069 & ~n0644;
assign n1449 =  n1447 & ~n1448;
assign n1450 =  n0055 & ~n0644;
assign n1451 =  n1449 & ~n1450;
assign n1452 =  n0054 & ~n0644;
assign n1453 =  n1451 & ~n1452;
assign n1454 =  n0053 & ~n0644;
assign n1455 =  n1453 & ~n1454;
assign n1456 =  n0052 & ~n0644;
assign n1457 =  n1455 & ~n1456;
assign n1458 =  n0049 & ~n0644;
assign n1459 =  n1457 & ~n1458;
assign n1460 =  n0391 & ~n0643;
assign n1461 =  n1459 & ~n1460;
assign n1462 =  n0407 & ~n0643;
assign n1463 =  n1461 & ~n1462;
assign n1464 =  n0392 & ~n0643;
assign n1465 =  n1463 & ~n1464;
assign n1466 =  n0393 & ~n0643;
assign n1467 =  n1465 & ~n1466;
assign n1468 =  n0394 & ~n0643;
assign n1469 =  n1467 & ~n1468;
assign n1470 =  n0408 & ~n0643;
assign n1471 =  n1469 & ~n1470;
assign n1472 =  n0409 & ~n0643;
assign n1473 =  n1471 & ~n1472;
assign n1474 =  n0410 & ~n0643;
assign n1475 =  n1473 & ~n1474;
assign n1476 =  n0072 & ~n0643;
assign n1477 =  n1475 & ~n1476;
assign n1478 =  n0066 & ~n0643;
assign n1479 =  n1477 & ~n1478;
assign n1480 =  n0042 & ~n0643;
assign n1481 =  n1479 & ~n1480;
assign n1482 =  n0041 & ~n0643;
assign n1483 =  n1481 & ~n1482;
assign n1484 =  n0040 & ~n0643;
assign n1485 =  n1483 & ~n1484;
assign n1486 =  n0039 & ~n0643;
assign n1487 =  n1485 & ~n1486;
assign n1488 =  n0036 & ~n0643;
assign n1489 =  n1487 & ~n1488;
assign n1490 =  n0386 & ~n0642;
assign n1491 =  n1489 & ~n1490;
assign n1492 =  n0387 & ~n0642;
assign n1493 =  n1491 & ~n1492;
assign n1494 =  n0402 & ~n0642;
assign n1495 =  n1493 & ~n1494;
assign n1496 =  n0403 & ~n0642;
assign n1497 =  n1495 & ~n1496;
assign n1498 =  n0388 & ~n0642;
assign n1499 =  n1497 & ~n1498;
assign n1500 =  n0404 & ~n0642;
assign n1501 =  n1499 & ~n1500;
assign n1502 =  n0389 & ~n0642;
assign n1503 =  n1501 & ~n1502;
assign n1504 =  n0405 & ~n0642;
assign n1505 =  n1503 & ~n1504;
assign n1506 =  n0071 & ~n0642;
assign n1507 =  n1505 & ~n1506;
assign n1508 =  n0063 & ~n0642;
assign n1509 =  n1507 & ~n1508;
assign n1510 =  n0029 & ~n0642;
assign n1511 =  n1509 & ~n1510;
assign n1512 =  n0028 & ~n0642;
assign n1513 =  n1511 & ~n1512;
assign n1514 =  n0027 & ~n0642;
assign n1515 =  n1513 & ~n1514;
assign n1516 =  n0026 & ~n0642;
assign n1517 =  n1515 & ~n1516;
assign n1518 =  n0023 & ~n0642;
assign n1519 =  n1517 & ~n1518;
assign n1520 =  n0640 &  n0898;
assign n1521 = ~n0641 &  n1520;
assign n1522 =  n1519 & ~n1521;
assign n1523 =  n0638 & ~n0640;
assign n1524 =  n1522 & ~n1523;
assign n1525 =  n0550 & ~n0640;
assign n1526 =  n1524 & ~n1525;
assign n1527 =  n0283 & ~n0640;
assign n1528 =  n1526 & ~n1527;
assign n1529 =  n0639 & ~n0640;
assign n1530 =  n1528 & ~n1529;
assign n1531 =  n0588 &  n0603;
assign n1532 = ~n0639 &  n1531;
assign n1533 =  n1530 & ~n1532;
assign n1534 =  n0637 &  n0912;
assign n1535 = ~n0638 &  n1534;
assign n1536 =  n1533 & ~n1535;
assign n1537 =  n0634 & ~n0637;
assign n1538 =  n1536 & ~n1537;
assign n1539 =  n0635 & ~n0637;
assign n1540 =  n1538 & ~n1539;
assign n1541 =  n0636 & ~n0637;
assign n1542 =  n1540 & ~n1541;
assign n1543 = ~n0069 &  n0924;
assign n1544 = ~n0049 &  n1543;
assign n1545 = ~n0073 &  n1544;
assign n1546 =  n0174 &  n1545;
assign n1547 =  n0190 &  n1546;
assign n1548 =  n0173 &  n1547;
assign n1549 =  n0189 &  n1548;
assign n1550 =  n0188 &  n1549;
assign n1551 =  n0172 &  n1550;
assign n1552 =  n0187 &  n1551;
assign n1553 =  n0171 &  n1552;
assign n1554 = ~n0636 &  n1553;
assign n1555 =  n1542 & ~n1554;
assign n1556 = ~n0036 & ~n0039;
assign n1557 = ~n0066 &  n1556;
assign n1558 = ~n0040 &  n1557;
assign n1559 = ~n0072 &  n1558;
assign n1560 = ~n0042 &  n1559;
assign n1561 = ~n0041 &  n1560;
assign n1562 =  n0185 &  n1561;
assign n1563 =  n0184 &  n1562;
assign n1564 =  n0183 &  n1563;
assign n1565 =  n0169 &  n1564;
assign n1566 =  n0168 &  n1565;
assign n1567 =  n0167 &  n1566;
assign n1568 =  n0182 &  n1567;
assign n1569 =  n0166 &  n1568;
assign n1570 = ~n0635 &  n1569;
assign n1571 =  n1555 & ~n1570;
assign n1572 = ~n0023 & ~n0028;
assign n1573 = ~n0029 &  n1572;
assign n1574 = ~n0027 &  n1573;
assign n1575 = ~n0026 &  n1574;
assign n1576 = ~n0063 &  n1575;
assign n1577 = ~n0071 &  n1576;
assign n1578 =  n0180 &  n1577;
assign n1579 =  n0164 &  n1578;
assign n1580 =  n0179 &  n1579;
assign n1581 =  n0163 &  n1580;
assign n1582 =  n0178 &  n1581;
assign n1583 =  n0177 &  n1582;
assign n1584 =  n0162 &  n1583;
assign n1585 =  n0161 &  n1584;
assign n1586 = ~n0634 &  n1585;
assign n1587 =  n1571 & ~n1586;
assign n1588 = ~n0002 &  n1025;
assign n1589 = ~n0001 &  n1588;
assign n1590 =  n0535 &  n1589;
assign n1591 =  n0534 &  n1590;
assign n1592 =  n0632 &  n1591;
assign n1593 = ~n0633 &  n1592;
assign n1594 =  n1587 & ~n1593;
assign n1595 =  n0628 & ~n0632;
assign n1596 =  n1594 & ~n1595;
assign n1597 =  n0631 & ~n0632;
assign n1598 =  n1596 & ~n1597;
assign n1599 =  n0478 &  n0531;
assign n1600 =  n0477 &  n1599;
assign n1601 =  n0476 &  n1600;
assign n1602 =  n0568 &  n1601;
assign n1603 =  n0566 &  n1602;
assign n1604 =  n0630 &  n1603;
assign n1605 =  n0629 &  n1604;
assign n1606 = ~n0631 &  n1605;
assign n1607 =  n1598 & ~n1606;
assign n1608 =  n0493 & ~n0630;
assign n1609 =  n1607 & ~n1608;
assign n1610 =  n0488 & ~n0630;
assign n1611 =  n1609 & ~n1610;
assign n1612 =  n0610 & ~n0629;
assign n1613 =  n1611 & ~n1612;
assign n1614 =  n0577 & ~n0629;
assign n1615 =  n1613 & ~n1614;
assign n1616 =  n0627 &  n0898;
assign n1617 = ~n0628 &  n1616;
assign n1618 =  n1615 & ~n1617;
assign n1619 =  n0625 & ~n0627;
assign n1620 =  n1618 & ~n1619;
assign n1621 =  n0626 & ~n0627;
assign n1622 =  n1620 & ~n1621;
assign n1623 =  n0542 & ~n0627;
assign n1624 =  n1622 & ~n1623;
assign n1625 =  n0544 & ~n0627;
assign n1626 =  n1624 & ~n1625;
assign n1627 =  n0251 & ~n0627;
assign n1628 =  n1626 & ~n1627;
assign n1629 =  n0252 & ~n0627;
assign n1630 =  n1628 & ~n1629;
assign n1631 =  n0253 & ~n0627;
assign n1632 =  n1630 & ~n1631;
assign n1633 =  n0263 &  n0268;
assign n1634 = ~n0626 &  n1633;
assign n1635 =  n1632 & ~n1634;
assign n1636 =  n0553 &  n0603;
assign n1637 = ~n0625 &  n1636;
assign n1638 =  n1635 & ~n1637;
assign n1639 = ~n0003 &  n1292;
assign n1640 = ~n0001 &  n1639;
assign n1641 =  n0535 &  n1640;
assign n1642 =  n0534 &  n1641;
assign n1643 =  n0623 &  n1642;
assign n1644 = ~n0624 &  n1643;
assign n1645 =  n1638 & ~n1644;
assign n1646 =  n0619 & ~n0623;
assign n1647 =  n1645 & ~n1646;
assign n1648 =  n0622 & ~n0623;
assign n1649 =  n1647 & ~n1648;
assign n1650 =  n0461 &  n0531;
assign n1651 =  n0460 &  n1650;
assign n1652 =  n0459 &  n1651;
assign n1653 =  n0458 &  n1652;
assign n1654 =  n0441 &  n1653;
assign n1655 =  n0621 &  n1654;
assign n1656 =  n0620 &  n1655;
assign n1657 = ~n0622 &  n1656;
assign n1658 =  n1649 & ~n1657;
assign n1659 =  n0493 & ~n0621;
assign n1660 =  n1658 & ~n1659;
assign n1661 =  n0573 & ~n0621;
assign n1662 =  n1660 & ~n1661;
assign n1663 =  n0581 & ~n0620;
assign n1664 =  n1662 & ~n1663;
assign n1665 =  n0511 & ~n0620;
assign n1666 =  n1664 & ~n1665;
assign n1667 =  n0618 &  n0898;
assign n1668 = ~n0619 &  n1667;
assign n1669 =  n1666 & ~n1668;
assign n1670 =  n0616 & ~n0618;
assign n1671 =  n1669 & ~n1670;
assign n1672 =  n0617 & ~n0618;
assign n1673 =  n1671 & ~n1672;
assign n1674 =  n0216 & ~n0618;
assign n1675 =  n1673 & ~n1674;
assign n1676 =  n0233 & ~n0618;
assign n1677 =  n1675 & ~n1676;
assign n1678 =  n0234 & ~n0618;
assign n1679 =  n1677 & ~n1678;
assign n1680 =  n0235 & ~n0618;
assign n1681 =  n1679 & ~n1680;
assign n1682 =  n0236 & ~n0618;
assign n1683 =  n1681 & ~n1682;
assign n1684 =  n0268 &  n0549;
assign n1685 = ~n0617 &  n1684;
assign n1686 =  n1683 & ~n1685;
assign n1687 =  n0286 &  n0557;
assign n1688 = ~n0616 &  n1687;
assign n1689 =  n1686 & ~n1688;
assign n1690 = ~n0001 &  n1080;
assign n1691 =  n0535 &  n1690;
assign n1692 =  n0534 &  n1691;
assign n1693 =  n0614 &  n1692;
assign n1694 = ~n0615 &  n1693;
assign n1695 =  n1689 & ~n1694;
assign n1696 =  n0607 & ~n0614;
assign n1697 =  n1695 & ~n1696;
assign n1698 =  n0613 & ~n0614;
assign n1699 =  n1697 & ~n1698;
assign n1700 =  n0516 &  n0531;
assign n1701 =  n0515 &  n1700;
assign n1702 =  n0514 &  n1701;
assign n1703 =  n0580 &  n1702;
assign n1704 =  n0579 &  n1703;
assign n1705 =  n0612 &  n1704;
assign n1706 =  n0611 &  n1705;
assign n1707 = ~n0613 &  n1706;
assign n1708 =  n1699 & ~n1707;
assign n1709 =  n0462 & ~n0612;
assign n1710 =  n1708 & ~n1709;
assign n1711 =  n0525 & ~n0612;
assign n1712 =  n1710 & ~n1711;
assign n1713 =  n0573 & ~n0611;
assign n1714 =  n1712 & ~n1713;
assign n1715 =  n0610 & ~n0611;
assign n1716 =  n1714 & ~n1715;
assign n1717 =  n0520 &  n0521;
assign n1718 =  n0519 &  n1717;
assign n1719 =  n0609 &  n1718;
assign n1720 =  n0608 &  n1719;
assign n1721 = ~n0610 &  n1720;
assign n1722 =  n1716 & ~n1721;
assign n1723 =  n0517 & ~n0609;
assign n1724 =  n1722 & ~n1723;
assign n1725 =  n0445 & ~n0609;
assign n1726 =  n1724 & ~n1725;
assign n1727 =  n0336 & ~n0609;
assign n1728 =  n1726 & ~n1727;
assign n1729 =  n0337 & ~n0609;
assign n1730 =  n1728 & ~n1729;
assign n1731 =  n0338 & ~n0609;
assign n1732 =  n1730 & ~n1731;
assign n1733 =  n0339 & ~n0609;
assign n1734 =  n1732 & ~n1733;
assign n1735 =  n0578 & ~n0608;
assign n1736 =  n1734 & ~n1735;
assign n1737 =  n0417 & ~n0608;
assign n1738 =  n1736 & ~n1737;
assign n1739 =  n0336 & ~n0608;
assign n1740 =  n1738 & ~n1739;
assign n1741 =  n0337 & ~n0608;
assign n1742 =  n1740 & ~n1741;
assign n1743 =  n0338 & ~n0608;
assign n1744 =  n1742 & ~n1743;
assign n1745 =  n0339 & ~n0608;
assign n1746 =  n1744 & ~n1745;
assign n1747 =  n0606 &  n0898;
assign n1748 = ~n0607 &  n1747;
assign n1749 =  n1746 & ~n1748;
assign n1750 =  n0604 & ~n0606;
assign n1751 =  n1749 & ~n1750;
assign n1752 =  n0605 & ~n0606;
assign n1753 =  n1751 & ~n1752;
assign n1754 =  n0555 & ~n0606;
assign n1755 =  n1753 & ~n1754;
assign n1756 =  n0556 & ~n0606;
assign n1757 =  n1755 & ~n1756;
assign n1758 =  n0289 & ~n0606;
assign n1759 =  n1757 & ~n1758;
assign n1760 =  n0290 & ~n0606;
assign n1761 =  n1759 & ~n1760;
assign n1762 =  n0291 & ~n0606;
assign n1763 =  n1761 & ~n1762;
assign n1764 =  n0237 &  n0300;
assign n1765 = ~n0605 &  n1764;
assign n1766 =  n1763 & ~n1765;
assign n1767 =  n0549 &  n0603;
assign n1768 = ~n0604 &  n1767;
assign n1769 =  n1766 & ~n1768;
assign n1770 =  n0601 & ~n0603;
assign n1771 =  n1769 & ~n1770;
assign n1772 =  n0602 & ~n0603;
assign n1773 =  n1771 & ~n1772;
assign n1774 =  n0294 & ~n0603;
assign n1775 =  n1773 & ~n1774;
assign n1776 =  n0295 & ~n0603;
assign n1777 =  n1775 & ~n1776;
assign n1778 =  n0296 & ~n0603;
assign n1779 =  n1777 & ~n1778;
assign n1780 =  n0220 &  n0912;
assign n1781 =  n0292 &  n1780;
assign n1782 = ~n0602 &  n1781;
assign n1783 =  n1779 & ~n1782;
assign n1784 =  n0192 &  n0912;
assign n1785 =  n0554 &  n1784;
assign n1786 = ~n0601 &  n1785;
assign n1787 =  n1783 & ~n1786;
assign n1788 = ~n0001 &  n1132;
assign n1789 =  n0535 &  n1788;
assign n1790 =  n0534 &  n1789;
assign n1791 =  n0599 &  n1790;
assign n1792 = ~n0600 &  n1791;
assign n1793 =  n1787 & ~n1792;
assign n1794 =  n0592 & ~n0599;
assign n1795 =  n1793 & ~n1794;
assign n1796 =  n0598 & ~n0599;
assign n1797 =  n1795 & ~n1796;
assign n1798 =  n0496 &  n0531;
assign n1799 =  n0495 &  n1798;
assign n1800 =  n0494 &  n1799;
assign n1801 =  n0572 &  n1800;
assign n1802 =  n0571 &  n1801;
assign n1803 =  n0597 &  n1802;
assign n1804 =  n0596 &  n1803;
assign n1805 = ~n0598 &  n1804;
assign n1806 =  n1797 & ~n1805;
assign n1807 =  n0462 & ~n0597;
assign n1808 =  n1806 & ~n1807;
assign n1809 =  n0507 & ~n0597;
assign n1810 =  n1808 & ~n1809;
assign n1811 =  n0595 & ~n0596;
assign n1812 =  n1810 & ~n1811;
assign n1813 =  n0581 & ~n0596;
assign n1814 =  n1812 & ~n1813;
assign n1815 =  n0501 &  n0594;
assign n1816 =  n0500 &  n1815;
assign n1817 =  n0499 &  n1816;
assign n1818 =  n0593 &  n1817;
assign n1819 = ~n0595 &  n1818;
assign n1820 =  n1814 & ~n1819;
assign n1821 =  n0497 & ~n0594;
assign n1822 =  n1820 & ~n1821;
assign n1823 =  n0368 & ~n0594;
assign n1824 =  n1822 & ~n1823;
assign n1825 =  n0336 & ~n0594;
assign n1826 =  n1824 & ~n1825;
assign n1827 =  n0337 & ~n0594;
assign n1828 =  n1826 & ~n1827;
assign n1829 =  n0338 & ~n0594;
assign n1830 =  n1828 & ~n1829;
assign n1831 =  n0339 & ~n0594;
assign n1832 =  n1830 & ~n1831;
assign n1833 =  n0570 & ~n0593;
assign n1834 =  n1832 & ~n1833;
assign n1835 =  n0422 & ~n0593;
assign n1836 =  n1834 & ~n1835;
assign n1837 =  n0336 & ~n0593;
assign n1838 =  n1836 & ~n1837;
assign n1839 =  n0337 & ~n0593;
assign n1840 =  n1838 & ~n1839;
assign n1841 =  n0338 & ~n0593;
assign n1842 =  n1840 & ~n1841;
assign n1843 =  n0339 & ~n0593;
assign n1844 =  n1842 & ~n1843;
assign n1845 =  n0591 &  n0898;
assign n1846 = ~n0592 &  n1845;
assign n1847 =  n1844 & ~n1846;
assign n1848 =  n0589 & ~n0591;
assign n1849 =  n1847 & ~n1848;
assign n1850 =  n0590 & ~n0591;
assign n1851 =  n1849 & ~n1850;
assign n1852 =  n0547 & ~n0591;
assign n1853 =  n1851 & ~n1852;
assign n1854 =  n0548 & ~n0591;
assign n1855 =  n1853 & ~n1854;
assign n1856 =  n0269 & ~n0591;
assign n1857 =  n1855 & ~n1856;
assign n1858 =  n0270 & ~n0591;
assign n1859 =  n1857 & ~n1858;
assign n1860 =  n0271 & ~n0591;
assign n1861 =  n1859 & ~n1860;
assign n1862 =  n0237 &  n0282;
assign n1863 = ~n0590 &  n1862;
assign n1864 =  n1861 & ~n1863;
assign n1865 =  n0557 &  n0588;
assign n1866 = ~n0589 &  n1865;
assign n1867 =  n1864 & ~n1866;
assign n1868 =  n0586 & ~n0588;
assign n1869 =  n1867 & ~n1868;
assign n1870 =  n0274 & ~n0588;
assign n1871 =  n1869 & ~n1870;
assign n1872 =  n0275 & ~n0588;
assign n1873 =  n1871 & ~n1872;
assign n1874 =  n0587 & ~n0588;
assign n1875 =  n1873 & ~n1874;
assign n1876 =  n0276 & ~n0588;
assign n1877 =  n1875 & ~n1876;
assign n1878 =  n0143 &  n0912;
assign n1879 =  n0272 &  n1878;
assign n1880 = ~n0587 &  n1879;
assign n1881 =  n1877 & ~n1880;
assign n1882 =  n0197 &  n0912;
assign n1883 =  n0546 &  n1882;
assign n1884 = ~n0586 &  n1883;
assign n1885 =  n1881 & ~n1884;
assign n1886 = ~n0001 &  n1026;
assign n1887 =  n0535 &  n1886;
assign n1888 =  n0534 &  n1887;
assign n1889 =  n0584 &  n1888;
assign n1890 = ~n0585 &  n1889;
assign n1891 =  n1885 & ~n1890;
assign n1892 =  n0560 & ~n0584;
assign n1893 =  n1891 & ~n1892;
assign n1894 =  n0583 & ~n0584;
assign n1895 =  n1893 & ~n1894;
assign n1896 =  n0531 &  n0582;
assign n1897 =  n0574 &  n1896;
assign n1898 =  n0489 &  n1897;
assign n1899 =  n0565 &  n1898;
assign n1900 = ~n0583 &  n1899;
assign n1901 =  n1895 & ~n1900;
assign n1902 =  n0577 & ~n0582;
assign n1903 =  n1901 & ~n1902;
assign n1904 =  n0581 & ~n0582;
assign n1905 =  n1903 & ~n1904;
assign n1906 =  n0515 &  n0516;
assign n1907 =  n0514 &  n1906;
assign n1908 =  n0580 &  n1907;
assign n1909 =  n0579 &  n1908;
assign n1910 = ~n0581 &  n1909;
assign n1911 =  n1905 & ~n1910;
assign n1912 =  n0457 & ~n0580;
assign n1913 =  n1911 & ~n1912;
assign n1914 =  n0522 & ~n0580;
assign n1915 =  n1913 & ~n1914;
assign n1916 =  n0336 & ~n0580;
assign n1917 =  n1915 & ~n1916;
assign n1918 =  n0337 & ~n0580;
assign n1919 =  n1917 & ~n1918;
assign n1920 =  n0338 & ~n0580;
assign n1921 =  n1919 & ~n1920;
assign n1922 =  n0339 & ~n0580;
assign n1923 =  n1921 & ~n1922;
assign n1924 =  n0578 & ~n0579;
assign n1925 =  n1923 & ~n1924;
assign n1926 =  n0384 & ~n0579;
assign n1927 =  n1925 & ~n1926;
assign n1928 =  n0336 & ~n0579;
assign n1929 =  n1927 & ~n1928;
assign n1930 =  n0337 & ~n0579;
assign n1931 =  n1929 & ~n1930;
assign n1932 =  n0338 & ~n0579;
assign n1933 =  n1931 & ~n1932;
assign n1934 =  n0339 & ~n0579;
assign n1935 =  n1933 & ~n1934;
assign n1936 =  n0513 &  n0524;
assign n1937 =  n0512 &  n1936;
assign n1938 = ~n0578 &  n1937;
assign n1939 =  n1935 & ~n1938;
assign n1940 =  n0469 &  n0576;
assign n1941 =  n0575 &  n1940;
assign n1942 =  n0468 &  n1941;
assign n1943 =  n0467 &  n1942;
assign n1944 = ~n0577 &  n1943;
assign n1945 =  n1939 & ~n1944;
assign n1946 =  n0479 & ~n0576;
assign n1947 =  n1945 & ~n1946;
assign n1948 =  n0401 & ~n0576;
assign n1949 =  n1947 & ~n1948;
assign n1950 =  n0336 & ~n0576;
assign n1951 =  n1949 & ~n1950;
assign n1952 =  n0337 & ~n0576;
assign n1953 =  n1951 & ~n1952;
assign n1954 =  n0338 & ~n0576;
assign n1955 =  n1953 & ~n1954;
assign n1956 =  n0339 & ~n0576;
assign n1957 =  n1955 & ~n1956;
assign n1958 =  n0567 & ~n0575;
assign n1959 =  n1957 & ~n1958;
assign n1960 =  n0422 & ~n0575;
assign n1961 =  n1959 & ~n1960;
assign n1962 =  n0336 & ~n0575;
assign n1963 =  n1961 & ~n1962;
assign n1964 =  n0337 & ~n0575;
assign n1965 =  n1963 & ~n1964;
assign n1966 =  n0338 & ~n0575;
assign n1967 =  n1965 & ~n1966;
assign n1968 =  n0339 & ~n0575;
assign n1969 =  n1967 & ~n1968;
assign n1970 =  n0569 & ~n0574;
assign n1971 =  n1969 & ~n1970;
assign n1972 =  n0573 & ~n0574;
assign n1973 =  n1971 & ~n1972;
assign n1974 =  n0495 &  n0496;
assign n1975 =  n0494 &  n1974;
assign n1976 =  n0572 &  n1975;
assign n1977 =  n0571 &  n1976;
assign n1978 = ~n0573 &  n1977;
assign n1979 =  n1973 & ~n1978;
assign n1980 =  n0502 & ~n0572;
assign n1981 =  n1979 & ~n1980;
assign n1982 =  n0440 & ~n0572;
assign n1983 =  n1981 & ~n1982;
assign n1984 =  n0336 & ~n0572;
assign n1985 =  n1983 & ~n1984;
assign n1986 =  n0337 & ~n0572;
assign n1987 =  n1985 & ~n1986;
assign n1988 =  n0338 & ~n0572;
assign n1989 =  n1987 & ~n1988;
assign n1990 =  n0339 & ~n0572;
assign n1991 =  n1989 & ~n1990;
assign n1992 =  n0570 & ~n0571;
assign n1993 =  n1991 & ~n1992;
assign n1994 =  n0384 & ~n0571;
assign n1995 =  n1993 & ~n1994;
assign n1996 =  n0336 & ~n0571;
assign n1997 =  n1995 & ~n1996;
assign n1998 =  n0337 & ~n0571;
assign n1999 =  n1997 & ~n1998;
assign n2000 =  n0338 & ~n0571;
assign n2001 =  n1999 & ~n2000;
assign n2002 =  n0339 & ~n0571;
assign n2003 =  n2001 & ~n2002;
assign n2004 =  n0505 &  n0506;
assign n2005 =  n0504 &  n2004;
assign n2006 = ~n0570 &  n2005;
assign n2007 =  n2003 & ~n2006;
assign n2008 =  n0477 &  n0478;
assign n2009 =  n0476 &  n2008;
assign n2010 =  n0568 &  n2009;
assign n2011 =  n0566 &  n2010;
assign n2012 = ~n0569 &  n2011;
assign n2013 =  n2007 & ~n2012;
assign n2014 =  n0567 & ~n0568;
assign n2015 =  n2013 & ~n2014;
assign n2016 =  n0417 & ~n0568;
assign n2017 =  n2015 & ~n2016;
assign n2018 =  n0336 & ~n0568;
assign n2019 =  n2017 & ~n2018;
assign n2020 =  n0337 & ~n0568;
assign n2021 =  n2019 & ~n2020;
assign n2022 =  n0338 & ~n0568;
assign n2023 =  n2021 & ~n2022;
assign n2024 =  n0339 & ~n0568;
assign n2025 =  n2023 & ~n2024;
assign n2026 =  n0486 &  n0487;
assign n2027 =  n0485 &  n2026;
assign n2028 = ~n0567 &  n2027;
assign n2029 =  n2025 & ~n2028;
assign n2030 =  n0470 & ~n0566;
assign n2031 =  n2029 & ~n2030;
assign n2032 =  n0450 & ~n0566;
assign n2033 =  n2031 & ~n2032;
assign n2034 =  n0336 & ~n0566;
assign n2035 =  n2033 & ~n2034;
assign n2036 =  n0337 & ~n0566;
assign n2037 =  n2035 & ~n2036;
assign n2038 =  n0338 & ~n0566;
assign n2039 =  n2037 & ~n2038;
assign n2040 =  n0339 & ~n0566;
assign n2041 =  n2039 & ~n2040;
assign n2042 =  n0564 & ~n0565;
assign n2043 =  n2041 & ~n2042;
assign n2044 =  n0336 & ~n0565;
assign n2045 =  n2043 & ~n2044;
assign n2046 =  n0337 & ~n0565;
assign n2047 =  n2045 & ~n2046;
assign n2048 =  n0338 & ~n0565;
assign n2049 =  n2047 & ~n2048;
assign n2050 =  n0339 & ~n0565;
assign n2051 =  n2049 & ~n2050;
assign n2052 =  n0562 &  n0563;
assign n2053 =  n0561 &  n2052;
assign n2054 = ~n0564 &  n2053;
assign n2055 =  n2051 & ~n2054;
assign n2056 =  n0379 & ~n0563;
assign n2057 =  n2055 & ~n2056;
assign n2058 =  n0360 & ~n0563;
assign n2059 =  n2057 & ~n2058;
assign n2060 =  n0361 & ~n0563;
assign n2061 =  n2059 & ~n2060;
assign n2062 =  n0364 & ~n0563;
assign n2063 =  n2061 & ~n2062;
assign n2064 =  n0366 & ~n0563;
assign n2065 =  n2063 & ~n2064;
assign n2066 =  n0380 & ~n0563;
assign n2067 =  n2065 & ~n2066;
assign n2068 =  n0381 & ~n0563;
assign n2069 =  n2067 & ~n2068;
assign n2070 =  n0073 & ~n0563;
assign n2071 =  n2069 & ~n2070;
assign n2072 =  n0069 & ~n0563;
assign n2073 =  n2071 & ~n2072;
assign n2074 =  n0055 & ~n0563;
assign n2075 =  n2073 & ~n2074;
assign n2076 =  n0054 & ~n0563;
assign n2077 =  n2075 & ~n2076;
assign n2078 =  n0053 & ~n0563;
assign n2079 =  n2077 & ~n2078;
assign n2080 =  n0052 & ~n0563;
assign n2081 =  n2079 & ~n2080;
assign n2082 =  n0049 & ~n0563;
assign n2083 =  n2081 & ~n2082;
assign n2084 =  n0382 & ~n0563;
assign n2085 =  n2083 & ~n2084;
assign n2086 =  n0350 & ~n0562;
assign n2087 =  n2085 & ~n2086;
assign n2088 =  n0351 & ~n0562;
assign n2089 =  n2087 & ~n2088;
assign n2090 =  n0353 & ~n0562;
assign n2091 =  n2089 & ~n2090;
assign n2092 =  n0355 & ~n0562;
assign n2093 =  n2091 & ~n2092;
assign n2094 =  n0374 & ~n0562;
assign n2095 =  n2093 & ~n2094;
assign n2096 =  n0375 & ~n0562;
assign n2097 =  n2095 & ~n2096;
assign n2098 =  n0376 & ~n0562;
assign n2099 =  n2097 & ~n2098;
assign n2100 =  n0072 & ~n0562;
assign n2101 =  n2099 & ~n2100;
assign n2102 =  n0066 & ~n0562;
assign n2103 =  n2101 & ~n2102;
assign n2104 =  n0042 & ~n0562;
assign n2105 =  n2103 & ~n2104;
assign n2106 =  n0041 & ~n0562;
assign n2107 =  n2105 & ~n2106;
assign n2108 =  n0040 & ~n0562;
assign n2109 =  n2107 & ~n2108;
assign n2110 =  n0377 & ~n0562;
assign n2111 =  n2109 & ~n2110;
assign n2112 =  n0039 & ~n0562;
assign n2113 =  n2111 & ~n2112;
assign n2114 =  n0036 & ~n0562;
assign n2115 =  n2113 & ~n2114;
assign n2116 =  n0342 & ~n0561;
assign n2117 =  n2115 & ~n2116;
assign n2118 =  n0343 & ~n0561;
assign n2119 =  n2117 & ~n2118;
assign n2120 =  n0344 & ~n0561;
assign n2121 =  n2119 & ~n2120;
assign n2122 =  n0369 & ~n0561;
assign n2123 =  n2121 & ~n2122;
assign n2124 =  n0370 & ~n0561;
assign n2125 =  n2123 & ~n2124;
assign n2126 =  n0371 & ~n0561;
assign n2127 =  n2125 & ~n2126;
assign n2128 =  n0347 & ~n0561;
assign n2129 =  n2127 & ~n2128;
assign n2130 =  n0372 & ~n0561;
assign n2131 =  n2129 & ~n2130;
assign n2132 =  n0071 & ~n0561;
assign n2133 =  n2131 & ~n2132;
assign n2134 =  n0063 & ~n0561;
assign n2135 =  n2133 & ~n2134;
assign n2136 =  n0029 & ~n0561;
assign n2137 =  n2135 & ~n2136;
assign n2138 =  n0028 & ~n0561;
assign n2139 =  n2137 & ~n2138;
assign n2140 =  n0027 & ~n0561;
assign n2141 =  n2139 & ~n2140;
assign n2142 =  n0026 & ~n0561;
assign n2143 =  n2141 & ~n2142;
assign n2144 =  n0023 & ~n0561;
assign n2145 =  n2143 & ~n2144;
assign n2146 =  n0559 &  n0898;
assign n2147 = ~n0560 &  n2146;
assign n2148 =  n2145 & ~n2147;
assign n2149 =  n0541 & ~n0559;
assign n2150 =  n2148 & ~n2149;
assign n2151 =  n0264 & ~n0559;
assign n2152 =  n2150 & ~n2151;
assign n2153 =  n0550 & ~n0559;
assign n2154 =  n2152 & ~n2153;
assign n2155 =  n0558 & ~n0559;
assign n2156 =  n2154 & ~n2155;
assign n2157 =  n0553 &  n0557;
assign n2158 = ~n0558 &  n2157;
assign n2159 =  n2156 & ~n2158;
assign n2160 =  n0555 & ~n0557;
assign n2161 =  n2159 & ~n2160;
assign n2162 =  n0556 & ~n0557;
assign n2163 =  n2161 & ~n2162;
assign n2164 =  n0289 & ~n0557;
assign n2165 =  n2163 & ~n2164;
assign n2166 =  n0290 & ~n0557;
assign n2167 =  n2165 & ~n2166;
assign n2168 =  n0291 & ~n0557;
assign n2169 =  n2167 & ~n2168;
assign n2170 =  n0297 &  n0912;
assign n2171 =  n0232 &  n2170;
assign n2172 = ~n0556 &  n2171;
assign n2173 =  n2169 & ~n2172;
assign n2174 =  n0159 &  n0912;
assign n2175 =  n0554 &  n2174;
assign n2176 = ~n0555 &  n2175;
assign n2177 =  n2173 & ~n2176;
assign n2178 =  n0287 & ~n0554;
assign n2179 =  n2177 & ~n2178;
assign n2180 =  n0288 & ~n0554;
assign n2181 =  n2179 & ~n2180;
assign n2182 =  n0299 & ~n0554;
assign n2183 =  n2181 & ~n2182;
assign n2184 =  n0242 & ~n0553;
assign n2185 =  n2183 & ~n2184;
assign n2186 =  n0243 & ~n0553;
assign n2187 =  n2185 & ~n2186;
assign n2188 =  n0551 & ~n0553;
assign n2189 =  n2187 & ~n2188;
assign n2190 =  n0552 & ~n0553;
assign n2191 =  n2189 & ~n2190;
assign n2192 =  n0244 & ~n0553;
assign n2193 =  n2191 & ~n2192;
assign n2194 =  n0176 &  n0912;
assign n2195 =  n0254 &  n2194;
assign n2196 = ~n0552 &  n2195;
assign n2197 =  n2193 & ~n2196;
assign n2198 =  n0543 &  n1882;
assign n2199 = ~n0551 &  n2198;
assign n2200 =  n2197 & ~n2199;
assign n2201 =  n0545 &  n0549;
assign n2202 = ~n0550 &  n2201;
assign n2203 =  n2200 & ~n2202;
assign n2204 =  n0547 & ~n0549;
assign n2205 =  n2203 & ~n2204;
assign n2206 =  n0548 & ~n0549;
assign n2207 =  n2205 & ~n2206;
assign n2208 =  n0269 & ~n0549;
assign n2209 =  n2207 & ~n2208;
assign n2210 =  n0270 & ~n0549;
assign n2211 =  n2209 & ~n2210;
assign n2212 =  n0271 & ~n0549;
assign n2213 =  n2211 & ~n2212;
assign n2214 =  n0215 &  n0912;
assign n2215 =  n0277 &  n2214;
assign n2216 = ~n0548 &  n2215;
assign n2217 =  n2213 & ~n2216;
assign n2218 =  n0546 &  n2174;
assign n2219 = ~n0547 &  n2218;
assign n2220 =  n2217 & ~n2219;
assign n2221 =  n0279 & ~n0546;
assign n2222 =  n2220 & ~n2221;
assign n2223 =  n0280 & ~n0546;
assign n2224 =  n2222 & ~n2223;
assign n2225 =  n0281 & ~n0546;
assign n2226 =  n2224 & ~n2225;
assign n2227 =  n0542 & ~n0545;
assign n2228 =  n2226 & ~n2227;
assign n2229 =  n0544 & ~n0545;
assign n2230 =  n2228 & ~n2229;
assign n2231 =  n0251 & ~n0545;
assign n2232 =  n2230 & ~n2231;
assign n2233 =  n0252 & ~n0545;
assign n2234 =  n2232 & ~n2233;
assign n2235 =  n0253 & ~n0545;
assign n2236 =  n2234 & ~n2235;
assign n2237 =  n0543 &  n1784;
assign n2238 = ~n0544 &  n2237;
assign n2239 =  n2236 & ~n2238;
assign n2240 =  n0260 & ~n0543;
assign n2241 =  n2239 & ~n2240;
assign n2242 =  n0261 & ~n0543;
assign n2243 =  n2241 & ~n2242;
assign n2244 =  n0262 & ~n0543;
assign n2245 =  n2243 & ~n2244;
assign n2246 =  n0225 &  n0912;
assign n2247 =  n0245 &  n2246;
assign n2248 = ~n0542 &  n2247;
assign n2249 =  n2245 & ~n2248;
assign n2250 =  n0540 &  n0912;
assign n2251 = ~n0541 &  n2250;
assign n2252 =  n2249 & ~n2251;
assign n2253 =  n0537 & ~n0540;
assign n2254 =  n2252 & ~n2253;
assign n2255 =  n0538 & ~n0540;
assign n2256 =  n2254 & ~n2255;
assign n2257 =  n0539 & ~n0540;
assign n2258 =  n2256 & ~n2257;
assign n2259 = ~n0054 &  n0157;
assign n2260 = ~n0053 &  n2259;
assign n2261 = ~n0055 &  n2260;
assign n2262 = ~n0052 &  n2261;
assign n2263 = ~n0069 &  n2262;
assign n2264 = ~n0049 &  n2263;
assign n2265 = ~n0073 &  n2264;
assign n2266 =  n0156 &  n2265;
assign n2267 =  n0155 &  n2266;
assign n2268 =  n0141 &  n2267;
assign n2269 =  n0139 &  n2268;
assign n2270 =  n0136 &  n2269;
assign n2271 =  n0135 &  n2270;
assign n2272 =  n0154 &  n2271;
assign n2273 = ~n0539 &  n2272;
assign n2274 =  n2258 & ~n2273;
assign n2275 = ~n0039 &  n0152;
assign n2276 = ~n0036 &  n2275;
assign n2277 = ~n0066 &  n2276;
assign n2278 = ~n0040 &  n2277;
assign n2279 = ~n0072 &  n2278;
assign n2280 = ~n0042 &  n2279;
assign n2281 = ~n0041 &  n2280;
assign n2282 =  n0151 &  n2281;
assign n2283 =  n0150 &  n2282;
assign n2284 =  n0149 &  n2283;
assign n2285 =  n0130 &  n2284;
assign n2286 =  n0128 &  n2285;
assign n2287 =  n0126 &  n2286;
assign n2288 =  n0125 &  n2287;
assign n2289 = ~n0538 &  n2288;
assign n2290 =  n2274 & ~n2289;
assign n2291 =  n0147 &  n1577;
assign n2292 =  n0146 &  n2291;
assign n2293 =  n0122 &  n2292;
assign n2294 =  n0145 &  n2293;
assign n2295 =  n0144 &  n2294;
assign n2296 =  n0119 &  n2295;
assign n2297 =  n0118 &  n2296;
assign n2298 =  n0117 &  n2297;
assign n2299 = ~n0537 &  n2298;
assign n2300 =  n2290 & ~n2299;
assign n2301 = ~n0002 &  n1639;
assign n2302 =  n0535 &  n2301;
assign n2303 =  n0534 &  n2302;
assign n2304 =  n0533 &  n2303;
assign n2305 = ~n0536 &  n2304;
assign n2306 =  n2300 & ~n2305;
assign n2307 =  n0007 & ~n0535;
assign n2308 =  n2306 & ~n2307;
assign n2309 =  n0003 & ~n0535;
assign n2310 =  n2308 & ~n2309;
assign n2311 =  n0002 & ~n0535;
assign n2312 =  n2310 & ~n2311;
assign n2313 =  n0001 & ~n0535;
assign n2314 =  n2312 & ~n2313;
assign n2315 =  n0008 & ~n0534;
assign n2316 =  n2314 & ~n2315;
assign n2317 =  n0006 & ~n0534;
assign n2318 =  n2316 & ~n2317;
assign n2319 =  n0005 & ~n0534;
assign n2320 =  n2318 & ~n2319;
assign n2321 =  n0004 & ~n0534;
assign n2322 =  n2320 & ~n2321;
assign n2323 =  n0307 & ~n0533;
assign n2324 =  n2322 & ~n2323;
assign n2325 =  n0532 & ~n0533;
assign n2326 =  n2324 & ~n2325;
assign n2327 =  n0508 &  n0786;
assign n2328 =  n0489 &  n2327;
assign n2329 =  n0340 &  n2328;
assign n2330 = ~n0532 &  n2329;
assign n2331 =  n2326 & ~n2330;
assign n2332 =  n0527 & ~n0531;
assign n2333 =  n2331 & ~n2332;
assign n2334 =  n0528 & ~n0531;
assign n2335 =  n2333 & ~n2334;
assign n2336 =  n0529 & ~n0531;
assign n2337 =  n2335 & ~n2336;
assign n2338 =  n0530 & ~n0531;
assign n2339 =  n2337 & ~n2338;
assign n2340 = ~n0013 & ~n0014;
assign n2341 = ~n0530 &  n2340;
assign n2342 =  n2339 & ~n2341;
assign n2343 = ~n0009 & ~n0010;
assign n2344 = ~n0529 &  n2343;
assign n2345 =  n2342 & ~n2344;
assign n2346 = ~n0011 & ~n0012;
assign n2347 = ~n0528 &  n2346;
assign n2348 =  n2345 & ~n2347;
assign n2349 = ~n0015 & ~n0016;
assign n2350 = ~n0527 &  n2349;
assign n2351 =  n2348 & ~n2350;
assign n2352 =  n0511 & ~n0526;
assign n2353 =  n2351 & ~n2352;
assign n2354 =  n0525 & ~n0526;
assign n2355 =  n2353 & ~n2354;
assign n2356 =  n0523 &  n0524;
assign n2357 =  n0518 &  n2356;
assign n2358 =  n0513 &  n2357;
assign n2359 =  n0512 &  n2358;
assign n2360 = ~n0525 &  n2359;
assign n2361 =  n2355 & ~n2360;
assign n2362 =  n0474 & ~n0524;
assign n2363 =  n2361 & ~n2362;
assign n2364 =  n0336 & ~n0524;
assign n2365 =  n2363 & ~n2364;
assign n2366 =  n0337 & ~n0524;
assign n2367 =  n2365 & ~n2366;
assign n2368 =  n0338 & ~n0524;
assign n2369 =  n2367 & ~n2368;
assign n2370 =  n0339 & ~n0524;
assign n2371 =  n2369 & ~n2370;
assign n2372 =  n0483 & ~n0523;
assign n2373 =  n2371 & ~n2372;
assign n2374 =  n0522 & ~n0523;
assign n2375 =  n2373 & ~n2374;
assign n2376 =  n0336 & ~n0523;
assign n2377 =  n2375 & ~n2376;
assign n2378 =  n0337 & ~n0523;
assign n2379 =  n2377 & ~n2378;
assign n2380 =  n0338 & ~n0523;
assign n2381 =  n2379 & ~n2380;
assign n2382 =  n0339 & ~n0523;
assign n2383 =  n2381 & ~n2382;
assign n2384 = ~n0522 &  n1718;
assign n2385 =  n2383 & ~n2384;
assign n2386 =  n0450 & ~n0521;
assign n2387 =  n2385 & ~n2386;
assign n2388 =  n0336 & ~n0521;
assign n2389 =  n2387 & ~n2388;
assign n2390 =  n0337 & ~n0521;
assign n2391 =  n2389 & ~n2390;
assign n2392 =  n0338 & ~n0521;
assign n2393 =  n2391 & ~n2392;
assign n2394 =  n0339 & ~n0521;
assign n2395 =  n2393 & ~n2394;
assign n2396 =  n0440 & ~n0520;
assign n2397 =  n2395 & ~n2396;
assign n2398 =  n0445 & ~n0520;
assign n2399 =  n2397 & ~n2398;
assign n2400 =  n0336 & ~n0520;
assign n2401 =  n2399 & ~n2400;
assign n2402 =  n0337 & ~n0520;
assign n2403 =  n2401 & ~n2402;
assign n2404 =  n0338 & ~n0520;
assign n2405 =  n2403 & ~n2404;
assign n2406 =  n0339 & ~n0520;
assign n2407 =  n2405 & ~n2406;
assign n2408 =  n0417 & ~n0519;
assign n2409 =  n2407 & ~n2408;
assign n2410 =  n0474 & ~n0519;
assign n2411 =  n2409 & ~n2410;
assign n2412 =  n0336 & ~n0519;
assign n2413 =  n2411 & ~n2412;
assign n2414 =  n0337 & ~n0519;
assign n2415 =  n2413 & ~n2414;
assign n2416 =  n0338 & ~n0519;
assign n2417 =  n2415 & ~n2416;
assign n2418 =  n0339 & ~n0519;
assign n2419 =  n2417 & ~n2418;
assign n2420 =  n0466 & ~n0518;
assign n2421 =  n2419 & ~n2420;
assign n2422 =  n0517 & ~n0518;
assign n2423 =  n2421 & ~n2422;
assign n2424 =  n0336 & ~n0518;
assign n2425 =  n2423 & ~n2424;
assign n2426 =  n0337 & ~n0518;
assign n2427 =  n2425 & ~n2426;
assign n2428 =  n0338 & ~n0518;
assign n2429 =  n2427 & ~n2428;
assign n2430 =  n0339 & ~n0518;
assign n2431 =  n2429 & ~n2430;
assign n2432 = ~n0517 &  n1907;
assign n2433 =  n2431 & ~n2432;
assign n2434 =  n0440 & ~n0516;
assign n2435 =  n2433 & ~n2434;
assign n2436 =  n0336 & ~n0516;
assign n2437 =  n2435 & ~n2436;
assign n2438 =  n0337 & ~n0516;
assign n2439 =  n2437 & ~n2438;
assign n2440 =  n0338 & ~n0516;
assign n2441 =  n2439 & ~n2440;
assign n2442 =  n0339 & ~n0516;
assign n2443 =  n2441 & ~n2442;
assign n2444 =  n0457 & ~n0515;
assign n2445 =  n2443 & ~n2444;
assign n2446 =  n0450 & ~n0515;
assign n2447 =  n2445 & ~n2446;
assign n2448 =  n0336 & ~n0515;
assign n2449 =  n2447 & ~n2448;
assign n2450 =  n0337 & ~n0515;
assign n2451 =  n2449 & ~n2450;
assign n2452 =  n0338 & ~n0515;
assign n2453 =  n2451 & ~n2452;
assign n2454 =  n0339 & ~n0515;
assign n2455 =  n2453 & ~n2454;
assign n2456 =  n0384 & ~n0514;
assign n2457 =  n2455 & ~n2456;
assign n2458 =  n0474 & ~n0514;
assign n2459 =  n2457 & ~n2458;
assign n2460 =  n0336 & ~n0514;
assign n2461 =  n2459 & ~n2460;
assign n2462 =  n0337 & ~n0514;
assign n2463 =  n2461 & ~n2462;
assign n2464 =  n0338 & ~n0514;
assign n2465 =  n2463 & ~n2464;
assign n2466 =  n0339 & ~n0514;
assign n2467 =  n2465 & ~n2466;
assign n2468 =  n0483 & ~n0513;
assign n2469 =  n2467 & ~n2468;
assign n2470 =  n0450 & ~n0513;
assign n2471 =  n2469 & ~n2470;
assign n2472 =  n0336 & ~n0513;
assign n2473 =  n2471 & ~n2472;
assign n2474 =  n0337 & ~n0513;
assign n2475 =  n2473 & ~n2474;
assign n2476 =  n0338 & ~n0513;
assign n2477 =  n2475 & ~n2476;
assign n2478 =  n0339 & ~n0513;
assign n2479 =  n2477 & ~n2478;
assign n2480 =  n0466 & ~n0512;
assign n2481 =  n2479 & ~n2480;
assign n2482 =  n0440 & ~n0512;
assign n2483 =  n2481 & ~n2482;
assign n2484 =  n0336 & ~n0512;
assign n2485 =  n2483 & ~n2484;
assign n2486 =  n0337 & ~n0512;
assign n2487 =  n2485 & ~n2486;
assign n2488 =  n0338 & ~n0512;
assign n2489 =  n2487 & ~n2488;
assign n2490 =  n0339 & ~n0512;
assign n2491 =  n2489 & ~n2490;
assign n2492 =  n0423 &  n0510;
assign n2493 =  n0509 &  n2492;
assign n2494 =  n0418 &  n2493;
assign n2495 =  n0385 &  n2494;
assign n2496 = ~n0511 &  n2495;
assign n2497 =  n2491 & ~n2496;
assign n2498 =  n0401 & ~n0510;
assign n2499 =  n2497 & ~n2498;
assign n2500 =  n0453 & ~n0510;
assign n2501 =  n2499 & ~n2500;
assign n2502 =  n0336 & ~n0510;
assign n2503 =  n2501 & ~n2502;
assign n2504 =  n0337 & ~n0510;
assign n2505 =  n2503 & ~n2504;
assign n2506 =  n0338 & ~n0510;
assign n2507 =  n2505 & ~n2506;
assign n2508 =  n0339 & ~n0510;
assign n2509 =  n2507 & ~n2508;
assign n2510 =  n0368 & ~n0509;
assign n2511 =  n2509 & ~n2510;
assign n2512 =  n0491 & ~n0509;
assign n2513 =  n2511 & ~n2512;
assign n2514 =  n0336 & ~n0509;
assign n2515 =  n2513 & ~n2514;
assign n2516 =  n0337 & ~n0509;
assign n2517 =  n2515 & ~n2516;
assign n2518 =  n0338 & ~n0509;
assign n2519 =  n2517 & ~n2518;
assign n2520 =  n0339 & ~n0509;
assign n2521 =  n2519 & ~n2520;
assign n2522 =  n0493 & ~n0508;
assign n2523 =  n2521 & ~n2522;
assign n2524 =  n0507 & ~n0508;
assign n2525 =  n2523 & ~n2524;
assign n2526 =  n0503 &  n2005;
assign n2527 =  n0498 &  n2526;
assign n2528 = ~n0507 &  n2527;
assign n2529 =  n2525 & ~n2528;
assign n2530 =  n0483 & ~n0506;
assign n2531 =  n2529 & ~n2530;
assign n2532 =  n0336 & ~n0506;
assign n2533 =  n2531 & ~n2532;
assign n2534 =  n0337 & ~n0506;
assign n2535 =  n2533 & ~n2534;
assign n2536 =  n0338 & ~n0506;
assign n2537 =  n2535 & ~n2536;
assign n2538 =  n0339 & ~n0506;
assign n2539 =  n2537 & ~n2538;
assign n2540 =  n0401 & ~n0505;
assign n2541 =  n2539 & ~n2540;
assign n2542 =  n0474 & ~n0505;
assign n2543 =  n2541 & ~n2542;
assign n2544 =  n0336 & ~n0505;
assign n2545 =  n2543 & ~n2544;
assign n2546 =  n0337 & ~n0505;
assign n2547 =  n2545 & ~n2546;
assign n2548 =  n0338 & ~n0505;
assign n2549 =  n2547 & ~n2548;
assign n2550 =  n0339 & ~n0505;
assign n2551 =  n2549 & ~n2550;
assign n2552 =  n0466 & ~n0504;
assign n2553 =  n2551 & ~n2552;
assign n2554 =  n0457 & ~n0504;
assign n2555 =  n2553 & ~n2554;
assign n2556 =  n0336 & ~n0504;
assign n2557 =  n2555 & ~n2556;
assign n2558 =  n0337 & ~n0504;
assign n2559 =  n2557 & ~n2558;
assign n2560 =  n0338 & ~n0504;
assign n2561 =  n2559 & ~n2560;
assign n2562 =  n0339 & ~n0504;
assign n2563 =  n2561 & ~n2562;
assign n2564 =  n0502 & ~n0503;
assign n2565 =  n2563 & ~n2564;
assign n2566 =  n0474 & ~n0503;
assign n2567 =  n2565 & ~n2566;
assign n2568 =  n0336 & ~n0503;
assign n2569 =  n2567 & ~n2568;
assign n2570 =  n0337 & ~n0503;
assign n2571 =  n2569 & ~n2570;
assign n2572 =  n0338 & ~n0503;
assign n2573 =  n2571 & ~n2572;
assign n2574 =  n0339 & ~n0503;
assign n2575 =  n2573 & ~n2574;
assign n2576 =  n0500 &  n0501;
assign n2577 =  n0499 &  n2576;
assign n2578 = ~n0502 &  n2577;
assign n2579 =  n2575 & ~n2578;
assign n2580 =  n0401 & ~n0501;
assign n2581 =  n2579 & ~n2580;
assign n2582 =  n0336 & ~n0501;
assign n2583 =  n2581 & ~n2582;
assign n2584 =  n0337 & ~n0501;
assign n2585 =  n2583 & ~n2584;
assign n2586 =  n0338 & ~n0501;
assign n2587 =  n2585 & ~n2586;
assign n2588 =  n0339 & ~n0501;
assign n2589 =  n2587 & ~n2588;
assign n2590 =  n0368 & ~n0500;
assign n2591 =  n2589 & ~n2590;
assign n2592 =  n0457 & ~n0500;
assign n2593 =  n2591 & ~n2592;
assign n2594 =  n0336 & ~n0500;
assign n2595 =  n2593 & ~n2594;
assign n2596 =  n0337 & ~n0500;
assign n2597 =  n2595 & ~n2596;
assign n2598 =  n0338 & ~n0500;
assign n2599 =  n2597 & ~n2598;
assign n2600 =  n0339 & ~n0500;
assign n2601 =  n2599 & ~n2600;
assign n2602 =  n0422 & ~n0499;
assign n2603 =  n2601 & ~n2602;
assign n2604 =  n0483 & ~n0499;
assign n2605 =  n2603 & ~n2604;
assign n2606 =  n0336 & ~n0499;
assign n2607 =  n2605 & ~n2606;
assign n2608 =  n0337 & ~n0499;
assign n2609 =  n2607 & ~n2608;
assign n2610 =  n0338 & ~n0499;
assign n2611 =  n2609 & ~n2610;
assign n2612 =  n0339 & ~n0499;
assign n2613 =  n2611 & ~n2612;
assign n2614 =  n0497 & ~n0498;
assign n2615 =  n2613 & ~n2614;
assign n2616 =  n0466 & ~n0498;
assign n2617 =  n2615 & ~n2616;
assign n2618 =  n0336 & ~n0498;
assign n2619 =  n2617 & ~n2618;
assign n2620 =  n0337 & ~n0498;
assign n2621 =  n2619 & ~n2620;
assign n2622 =  n0338 & ~n0498;
assign n2623 =  n2621 & ~n2622;
assign n2624 =  n0339 & ~n0498;
assign n2625 =  n2623 & ~n2624;
assign n2626 = ~n0497 &  n1975;
assign n2627 =  n2625 & ~n2626;
assign n2628 =  n0457 & ~n0496;
assign n2629 =  n2627 & ~n2628;
assign n2630 =  n0336 & ~n0496;
assign n2631 =  n2629 & ~n2630;
assign n2632 =  n0337 & ~n0496;
assign n2633 =  n2631 & ~n2632;
assign n2634 =  n0338 & ~n0496;
assign n2635 =  n2633 & ~n2634;
assign n2636 =  n0339 & ~n0496;
assign n2637 =  n2635 & ~n2636;
assign n2638 =  n0401 & ~n0495;
assign n2639 =  n2637 & ~n2638;
assign n2640 =  n0440 & ~n0495;
assign n2641 =  n2639 & ~n2640;
assign n2642 =  n0336 & ~n0495;
assign n2643 =  n2641 & ~n2642;
assign n2644 =  n0337 & ~n0495;
assign n2645 =  n2643 & ~n2644;
assign n2646 =  n0338 & ~n0495;
assign n2647 =  n2645 & ~n2646;
assign n2648 =  n0339 & ~n0495;
assign n2649 =  n2647 & ~n2648;
assign n2650 =  n0384 & ~n0494;
assign n2651 =  n2649 & ~n2650;
assign n2652 =  n0483 & ~n0494;
assign n2653 =  n2651 & ~n2652;
assign n2654 =  n0336 & ~n0494;
assign n2655 =  n2653 & ~n2654;
assign n2656 =  n0337 & ~n0494;
assign n2657 =  n2655 & ~n2656;
assign n2658 =  n0338 & ~n0494;
assign n2659 =  n2657 & ~n2658;
assign n2660 =  n0339 & ~n0494;
assign n2661 =  n2659 & ~n2660;
assign n2662 =  n0451 &  n0452;
assign n2663 =  n0446 &  n2662;
assign n2664 =  n0492 &  n2663;
assign n2665 =  n0490 &  n2664;
assign n2666 = ~n0493 &  n2665;
assign n2667 =  n2661 & ~n2666;
assign n2668 =  n0491 & ~n0492;
assign n2669 =  n2667 & ~n2668;
assign n2670 =  n0445 & ~n0492;
assign n2671 =  n2669 & ~n2670;
assign n2672 =  n0336 & ~n0492;
assign n2673 =  n2671 & ~n2672;
assign n2674 =  n0337 & ~n0492;
assign n2675 =  n2673 & ~n2674;
assign n2676 =  n0338 & ~n0492;
assign n2677 =  n2675 & ~n2676;
assign n2678 =  n0339 & ~n0492;
assign n2679 =  n2677 & ~n2678;
assign n2680 =  n0460 &  n0461;
assign n2681 =  n0459 &  n2680;
assign n2682 = ~n0491 &  n2681;
assign n2683 =  n2679 & ~n2682;
assign n2684 =  n0424 & ~n0490;
assign n2685 =  n2683 & ~n2684;
assign n2686 =  n0450 & ~n0490;
assign n2687 =  n2685 & ~n2686;
assign n2688 =  n0336 & ~n0490;
assign n2689 =  n2687 & ~n2688;
assign n2690 =  n0337 & ~n0490;
assign n2691 =  n2689 & ~n2690;
assign n2692 =  n0338 & ~n0490;
assign n2693 =  n2691 & ~n2692;
assign n2694 =  n0339 & ~n0490;
assign n2695 =  n2693 & ~n2694;
assign n2696 =  n0462 & ~n0489;
assign n2697 =  n2695 & ~n2696;
assign n2698 =  n0488 & ~n0489;
assign n2699 =  n2697 & ~n2698;
assign n2700 =  n0484 &  n2027;
assign n2701 =  n0475 &  n2700;
assign n2702 = ~n0488 &  n2701;
assign n2703 =  n2699 & ~n2702;
assign n2704 =  n0466 & ~n0487;
assign n2705 =  n2703 & ~n2704;
assign n2706 =  n0336 & ~n0487;
assign n2707 =  n2705 & ~n2706;
assign n2708 =  n0337 & ~n0487;
assign n2709 =  n2707 & ~n2708;
assign n2710 =  n0338 & ~n0487;
assign n2711 =  n2709 & ~n2710;
assign n2712 =  n0339 & ~n0487;
assign n2713 =  n2711 & ~n2712;
assign n2714 =  n0368 & ~n0486;
assign n2715 =  n2713 & ~n2714;
assign n2716 =  n0474 & ~n0486;
assign n2717 =  n2715 & ~n2716;
assign n2718 =  n0336 & ~n0486;
assign n2719 =  n2717 & ~n2718;
assign n2720 =  n0337 & ~n0486;
assign n2721 =  n2719 & ~n2720;
assign n2722 =  n0338 & ~n0486;
assign n2723 =  n2721 & ~n2722;
assign n2724 =  n0339 & ~n0486;
assign n2725 =  n2723 & ~n2724;
assign n2726 =  n0483 & ~n0485;
assign n2727 =  n2725 & ~n2726;
assign n2728 =  n0445 & ~n0485;
assign n2729 =  n2727 & ~n2728;
assign n2730 =  n0336 & ~n0485;
assign n2731 =  n2729 & ~n2730;
assign n2732 =  n0337 & ~n0485;
assign n2733 =  n2731 & ~n2732;
assign n2734 =  n0338 & ~n0485;
assign n2735 =  n2733 & ~n2734;
assign n2736 =  n0339 & ~n0485;
assign n2737 =  n2735 & ~n2736;
assign n2738 =  n0479 & ~n0484;
assign n2739 =  n2737 & ~n2738;
assign n2740 =  n0483 & ~n0484;
assign n2741 =  n2739 & ~n2740;
assign n2742 =  n0336 & ~n0484;
assign n2743 =  n2741 & ~n2742;
assign n2744 =  n0337 & ~n0484;
assign n2745 =  n2743 & ~n2744;
assign n2746 =  n0338 & ~n0484;
assign n2747 =  n2745 & ~n2746;
assign n2748 =  n0339 & ~n0484;
assign n2749 =  n2747 & ~n2748;
assign n2750 =  n0481 &  n0482;
assign n2751 =  n0480 &  n2750;
assign n2752 = ~n0483 &  n2751;
assign n2753 =  n2749 & ~n2752;
assign n2754 =  n0396 & ~n0482;
assign n2755 =  n2753 & ~n2754;
assign n2756 =  n0328 & ~n0482;
assign n2757 =  n2755 & ~n2756;
assign n2758 =  n0330 & ~n0482;
assign n2759 =  n2757 & ~n2758;
assign n2760 =  n0331 & ~n0482;
assign n2761 =  n2759 & ~n2760;
assign n2762 =  n0397 & ~n0482;
assign n2763 =  n2761 & ~n2762;
assign n2764 =  n0332 & ~n0482;
assign n2765 =  n2763 & ~n2764;
assign n2766 =  n0398 & ~n0482;
assign n2767 =  n2765 & ~n2766;
assign n2768 =  n0399 & ~n0482;
assign n2769 =  n2767 & ~n2768;
assign n2770 =  n0082 & ~n0482;
assign n2771 =  n2769 & ~n2770;
assign n2772 =  n0073 & ~n0482;
assign n2773 =  n2771 & ~n2772;
assign n2774 =  n0069 & ~n0482;
assign n2775 =  n2773 & ~n2774;
assign n2776 =  n0068 & ~n0482;
assign n2777 =  n2775 & ~n2776;
assign n2778 =  n0055 & ~n0482;
assign n2779 =  n2777 & ~n2778;
assign n2780 =  n0054 & ~n0482;
assign n2781 =  n2779 & ~n2780;
assign n2782 =  n0053 & ~n0482;
assign n2783 =  n2781 & ~n2782;
assign n2784 =  n0391 & ~n0481;
assign n2785 =  n2783 & ~n2784;
assign n2786 =  n0319 & ~n0481;
assign n2787 =  n2785 & ~n2786;
assign n2788 =  n0320 & ~n0481;
assign n2789 =  n2787 & ~n2788;
assign n2790 =  n0392 & ~n0481;
assign n2791 =  n2789 & ~n2790;
assign n2792 =  n0393 & ~n0481;
assign n2793 =  n2791 & ~n2792;
assign n2794 =  n0394 & ~n0481;
assign n2795 =  n2793 & ~n2794;
assign n2796 =  n0322 & ~n0481;
assign n2797 =  n2795 & ~n2796;
assign n2798 =  n0324 & ~n0481;
assign n2799 =  n2797 & ~n2798;
assign n2800 =  n0081 & ~n0481;
assign n2801 =  n2799 & ~n2800;
assign n2802 =  n0072 & ~n0481;
assign n2803 =  n2801 & ~n2802;
assign n2804 =  n0066 & ~n0481;
assign n2805 =  n2803 & ~n2804;
assign n2806 =  n0065 & ~n0481;
assign n2807 =  n2805 & ~n2806;
assign n2808 =  n0042 & ~n0481;
assign n2809 =  n2807 & ~n2808;
assign n2810 =  n0041 & ~n0481;
assign n2811 =  n2809 & ~n2810;
assign n2812 =  n0040 & ~n0481;
assign n2813 =  n2811 & ~n2812;
assign n2814 =  n0386 & ~n0480;
assign n2815 =  n2813 & ~n2814;
assign n2816 =  n0387 & ~n0480;
assign n2817 =  n2815 & ~n2816;
assign n2818 =  n0309 & ~n0480;
assign n2819 =  n2817 & ~n2818;
assign n2820 =  n0310 & ~n0480;
assign n2821 =  n2819 & ~n2820;
assign n2822 =  n0313 & ~n0480;
assign n2823 =  n2821 & ~n2822;
assign n2824 =  n0388 & ~n0480;
assign n2825 =  n2823 & ~n2824;
assign n2826 =  n0389 & ~n0480;
assign n2827 =  n2825 & ~n2826;
assign n2828 =  n0314 & ~n0480;
assign n2829 =  n2827 & ~n2828;
assign n2830 =  n0080 & ~n0480;
assign n2831 =  n2829 & ~n2830;
assign n2832 =  n0071 & ~n0480;
assign n2833 =  n2831 & ~n2832;
assign n2834 =  n0063 & ~n0480;
assign n2835 =  n2833 & ~n2834;
assign n2836 =  n0062 & ~n0480;
assign n2837 =  n2835 & ~n2836;
assign n2838 =  n0029 & ~n0480;
assign n2839 =  n2837 & ~n2838;
assign n2840 =  n0028 & ~n0480;
assign n2841 =  n2839 & ~n2840;
assign n2842 =  n0027 & ~n0480;
assign n2843 =  n2841 & ~n2842;
assign n2844 = ~n0479 &  n2009;
assign n2845 =  n2843 & ~n2844;
assign n2846 =  n0445 & ~n0478;
assign n2847 =  n2845 & ~n2846;
assign n2848 =  n0336 & ~n0478;
assign n2849 =  n2847 & ~n2848;
assign n2850 =  n0337 & ~n0478;
assign n2851 =  n2849 & ~n2850;
assign n2852 =  n0338 & ~n0478;
assign n2853 =  n2851 & ~n2852;
assign n2854 =  n0339 & ~n0478;
assign n2855 =  n2853 & ~n2854;
assign n2856 =  n0368 & ~n0477;
assign n2857 =  n2855 & ~n2856;
assign n2858 =  n0450 & ~n0477;
assign n2859 =  n2857 & ~n2858;
assign n2860 =  n0336 & ~n0477;
assign n2861 =  n2859 & ~n2860;
assign n2862 =  n0337 & ~n0477;
assign n2863 =  n2861 & ~n2862;
assign n2864 =  n0338 & ~n0477;
assign n2865 =  n2863 & ~n2864;
assign n2866 =  n0339 & ~n0477;
assign n2867 =  n2865 & ~n2866;
assign n2868 =  n0466 & ~n0476;
assign n2869 =  n2867 & ~n2868;
assign n2870 =  n0417 & ~n0476;
assign n2871 =  n2869 & ~n2870;
assign n2872 =  n0336 & ~n0476;
assign n2873 =  n2871 & ~n2872;
assign n2874 =  n0337 & ~n0476;
assign n2875 =  n2873 & ~n2874;
assign n2876 =  n0338 & ~n0476;
assign n2877 =  n2875 & ~n2876;
assign n2878 =  n0339 & ~n0476;
assign n2879 =  n2877 & ~n2878;
assign n2880 =  n0470 & ~n0475;
assign n2881 =  n2879 & ~n2880;
assign n2882 =  n0474 & ~n0475;
assign n2883 =  n2881 & ~n2882;
assign n2884 =  n0336 & ~n0475;
assign n2885 =  n2883 & ~n2884;
assign n2886 =  n0337 & ~n0475;
assign n2887 =  n2885 & ~n2886;
assign n2888 =  n0338 & ~n0475;
assign n2889 =  n2887 & ~n2888;
assign n2890 =  n0339 & ~n0475;
assign n2891 =  n2889 & ~n2890;
assign n2892 =  n0472 &  n0473;
assign n2893 =  n0471 &  n2892;
assign n2894 = ~n0474 &  n2893;
assign n2895 =  n2891 & ~n2894;
assign n2896 =  n0435 & ~n0473;
assign n2897 =  n2895 & ~n2896;
assign n2898 =  n0328 & ~n0473;
assign n2899 =  n2897 & ~n2898;
assign n2900 =  n0330 & ~n0473;
assign n2901 =  n2899 & ~n2900;
assign n2902 =  n0331 & ~n0473;
assign n2903 =  n2901 & ~n2902;
assign n2904 =  n0436 & ~n0473;
assign n2905 =  n2903 & ~n2904;
assign n2906 =  n0332 & ~n0473;
assign n2907 =  n2905 & ~n2906;
assign n2908 =  n0437 & ~n0473;
assign n2909 =  n2907 & ~n2908;
assign n2910 =  n0438 & ~n0473;
assign n2911 =  n2909 & ~n2910;
assign n2912 =  n0082 & ~n0473;
assign n2913 =  n2911 & ~n2912;
assign n2914 =  n0073 & ~n0473;
assign n2915 =  n2913 & ~n2914;
assign n2916 =  n0068 & ~n0473;
assign n2917 =  n2915 & ~n2916;
assign n2918 =  n0055 & ~n0473;
assign n2919 =  n2917 & ~n2918;
assign n2920 =  n0054 & ~n0473;
assign n2921 =  n2919 & ~n2920;
assign n2922 =  n0053 & ~n0473;
assign n2923 =  n2921 & ~n2922;
assign n2924 =  n0051 & ~n0473;
assign n2925 =  n2923 & ~n2924;
assign n2926 =  n0430 & ~n0472;
assign n2927 =  n2925 & ~n2926;
assign n2928 =  n0431 & ~n0472;
assign n2929 =  n2927 & ~n2928;
assign n2930 =  n0432 & ~n0472;
assign n2931 =  n2929 & ~n2930;
assign n2932 =  n0319 & ~n0472;
assign n2933 =  n2931 & ~n2932;
assign n2934 =  n0320 & ~n0472;
assign n2935 =  n2933 & ~n2934;
assign n2936 =  n0433 & ~n0472;
assign n2937 =  n2935 & ~n2936;
assign n2938 =  n0322 & ~n0472;
assign n2939 =  n2937 & ~n2938;
assign n2940 =  n0324 & ~n0472;
assign n2941 =  n2939 & ~n2940;
assign n2942 =  n0081 & ~n0472;
assign n2943 =  n2941 & ~n2942;
assign n2944 =  n0072 & ~n0472;
assign n2945 =  n2943 & ~n2944;
assign n2946 =  n0065 & ~n0472;
assign n2947 =  n2945 & ~n2946;
assign n2948 =  n0042 & ~n0472;
assign n2949 =  n2947 & ~n2948;
assign n2950 =  n0041 & ~n0472;
assign n2951 =  n2949 & ~n2950;
assign n2952 =  n0040 & ~n0472;
assign n2953 =  n2951 & ~n2952;
assign n2954 =  n0038 & ~n0472;
assign n2955 =  n2953 & ~n2954;
assign n2956 =  n0425 & ~n0471;
assign n2957 =  n2955 & ~n2956;
assign n2958 =  n0426 & ~n0471;
assign n2959 =  n2957 & ~n2958;
assign n2960 =  n0427 & ~n0471;
assign n2961 =  n2959 & ~n2960;
assign n2962 =  n0309 & ~n0471;
assign n2963 =  n2961 & ~n2962;
assign n2964 =  n0310 & ~n0471;
assign n2965 =  n2963 & ~n2964;
assign n2966 =  n0313 & ~n0471;
assign n2967 =  n2965 & ~n2966;
assign n2968 =  n0314 & ~n0471;
assign n2969 =  n2967 & ~n2968;
assign n2970 =  n0080 & ~n0471;
assign n2971 =  n2969 & ~n2970;
assign n2972 =  n0071 & ~n0471;
assign n2973 =  n2971 & ~n2972;
assign n2974 =  n0062 & ~n0471;
assign n2975 =  n2973 & ~n2974;
assign n2976 =  n0428 & ~n0471;
assign n2977 =  n2975 & ~n2976;
assign n2978 =  n0029 & ~n0471;
assign n2979 =  n2977 & ~n2978;
assign n2980 =  n0028 & ~n0471;
assign n2981 =  n2979 & ~n2980;
assign n2982 =  n0027 & ~n0471;
assign n2983 =  n2981 & ~n2982;
assign n2984 =  n0025 & ~n0471;
assign n2985 =  n2983 & ~n2984;
assign n2986 =  n0468 &  n0469;
assign n2987 =  n0467 &  n2986;
assign n2988 = ~n0470 &  n2987;
assign n2989 =  n2985 & ~n2988;
assign n2990 =  n0368 & ~n0469;
assign n2991 =  n2989 & ~n2990;
assign n2992 =  n0336 & ~n0469;
assign n2993 =  n2991 & ~n2992;
assign n2994 =  n0337 & ~n0469;
assign n2995 =  n2993 & ~n2994;
assign n2996 =  n0338 & ~n0469;
assign n2997 =  n2995 & ~n2996;
assign n2998 =  n0339 & ~n0469;
assign n2999 =  n2997 & ~n2998;
assign n3000 =  n0401 & ~n0468;
assign n3001 =  n2999 & ~n3000;
assign n3002 =  n0445 & ~n0468;
assign n3003 =  n3001 & ~n3002;
assign n3004 =  n0336 & ~n0468;
assign n3005 =  n3003 & ~n3004;
assign n3006 =  n0337 & ~n0468;
assign n3007 =  n3005 & ~n3006;
assign n3008 =  n0338 & ~n0468;
assign n3009 =  n3007 & ~n3008;
assign n3010 =  n0339 & ~n0468;
assign n3011 =  n3009 & ~n3010;
assign n3012 =  n0422 & ~n0467;
assign n3013 =  n3011 & ~n3012;
assign n3014 =  n0466 & ~n0467;
assign n3015 =  n3013 & ~n3014;
assign n3016 =  n0336 & ~n0467;
assign n3017 =  n3015 & ~n3016;
assign n3018 =  n0337 & ~n0467;
assign n3019 =  n3017 & ~n3018;
assign n3020 =  n0338 & ~n0467;
assign n3021 =  n3019 & ~n3020;
assign n3022 =  n0339 & ~n0467;
assign n3023 =  n3021 & ~n3022;
assign n3024 =  n0464 &  n0465;
assign n3025 =  n0463 &  n3024;
assign n3026 = ~n0466 &  n3025;
assign n3027 =  n3023 & ~n3026;
assign n3028 =  n0360 & ~n0465;
assign n3029 =  n3027 & ~n3028;
assign n3030 =  n0361 & ~n0465;
assign n3031 =  n3029 & ~n3030;
assign n3032 =  n0364 & ~n0465;
assign n3033 =  n3031 & ~n3032;
assign n3034 =  n0328 & ~n0465;
assign n3035 =  n3033 & ~n3034;
assign n3036 =  n0330 & ~n0465;
assign n3037 =  n3035 & ~n3036;
assign n3038 =  n0331 & ~n0465;
assign n3039 =  n3037 & ~n3038;
assign n3040 =  n0366 & ~n0465;
assign n3041 =  n3039 & ~n3040;
assign n3042 =  n0332 & ~n0465;
assign n3043 =  n3041 & ~n3042;
assign n3044 =  n0082 & ~n0465;
assign n3045 =  n3043 & ~n3044;
assign n3046 =  n0076 & ~n0465;
assign n3047 =  n3045 & ~n3046;
assign n3048 =  n0073 & ~n0465;
assign n3049 =  n3047 & ~n3048;
assign n3050 =  n0069 & ~n0465;
assign n3051 =  n3049 & ~n3050;
assign n3052 =  n0068 & ~n0465;
assign n3053 =  n3051 & ~n3052;
assign n3054 =  n0054 & ~n0465;
assign n3055 =  n3053 & ~n3054;
assign n3056 =  n0053 & ~n0465;
assign n3057 =  n3055 & ~n3056;
assign n3058 =  n0350 & ~n0464;
assign n3059 =  n3057 & ~n3058;
assign n3060 =  n0351 & ~n0464;
assign n3061 =  n3059 & ~n3060;
assign n3062 =  n0353 & ~n0464;
assign n3063 =  n3061 & ~n3062;
assign n3064 =  n0355 & ~n0464;
assign n3065 =  n3063 & ~n3064;
assign n3066 =  n0319 & ~n0464;
assign n3067 =  n3065 & ~n3066;
assign n3068 =  n0320 & ~n0464;
assign n3069 =  n3067 & ~n3068;
assign n3070 =  n0322 & ~n0464;
assign n3071 =  n3069 & ~n3070;
assign n3072 =  n0324 & ~n0464;
assign n3073 =  n3071 & ~n3072;
assign n3074 =  n0081 & ~n0464;
assign n3075 =  n3073 & ~n3074;
assign n3076 =  n0075 & ~n0464;
assign n3077 =  n3075 & ~n3076;
assign n3078 =  n0072 & ~n0464;
assign n3079 =  n3077 & ~n3078;
assign n3080 =  n0066 & ~n0464;
assign n3081 =  n3079 & ~n3080;
assign n3082 =  n0065 & ~n0464;
assign n3083 =  n3081 & ~n3082;
assign n3084 =  n0041 & ~n0464;
assign n3085 =  n3083 & ~n3084;
assign n3086 =  n0040 & ~n0464;
assign n3087 =  n3085 & ~n3086;
assign n3088 =  n0342 & ~n0463;
assign n3089 =  n3087 & ~n3088;
assign n3090 =  n0343 & ~n0463;
assign n3091 =  n3089 & ~n3090;
assign n3092 =  n0344 & ~n0463;
assign n3093 =  n3091 & ~n3092;
assign n3094 =  n0309 & ~n0463;
assign n3095 =  n3093 & ~n3094;
assign n3096 =  n0310 & ~n0463;
assign n3097 =  n3095 & ~n3096;
assign n3098 =  n0313 & ~n0463;
assign n3099 =  n3097 & ~n3098;
assign n3100 =  n0347 & ~n0463;
assign n3101 =  n3099 & ~n3100;
assign n3102 =  n0314 & ~n0463;
assign n3103 =  n3101 & ~n3102;
assign n3104 =  n0080 & ~n0463;
assign n3105 =  n3103 & ~n3104;
assign n3106 =  n0074 & ~n0463;
assign n3107 =  n3105 & ~n3106;
assign n3108 =  n0071 & ~n0463;
assign n3109 =  n3107 & ~n3108;
assign n3110 =  n0063 & ~n0463;
assign n3111 =  n3109 & ~n3110;
assign n3112 =  n0062 & ~n0463;
assign n3113 =  n3111 & ~n3112;
assign n3114 =  n0028 & ~n0463;
assign n3115 =  n3113 & ~n3114;
assign n3116 =  n0027 & ~n0463;
assign n3117 =  n3115 & ~n3116;
assign n3118 =  n0458 &  n2681;
assign n3119 =  n0441 &  n3118;
assign n3120 = ~n0462 &  n3119;
assign n3121 =  n3117 & ~n3120;
assign n3122 =  n0384 & ~n0461;
assign n3123 =  n3121 & ~n3122;
assign n3124 =  n0336 & ~n0461;
assign n3125 =  n3123 & ~n3124;
assign n3126 =  n0337 & ~n0461;
assign n3127 =  n3125 & ~n3126;
assign n3128 =  n0338 & ~n0461;
assign n3129 =  n3127 & ~n3128;
assign n3130 =  n0339 & ~n0461;
assign n3131 =  n3129 & ~n3130;
assign n3132 =  n0422 & ~n0460;
assign n3133 =  n3131 & ~n3132;
assign n3134 =  n0440 & ~n0460;
assign n3135 =  n3133 & ~n3134;
assign n3136 =  n0336 & ~n0460;
assign n3137 =  n3135 & ~n3136;
assign n3138 =  n0337 & ~n0460;
assign n3139 =  n3137 & ~n3138;
assign n3140 =  n0338 & ~n0460;
assign n3141 =  n3139 & ~n3140;
assign n3142 =  n0339 & ~n0460;
assign n3143 =  n3141 & ~n3142;
assign n3144 =  n0457 & ~n0459;
assign n3145 =  n3143 & ~n3144;
assign n3146 =  n0417 & ~n0459;
assign n3147 =  n3145 & ~n3146;
assign n3148 =  n0336 & ~n0459;
assign n3149 =  n3147 & ~n3148;
assign n3150 =  n0337 & ~n0459;
assign n3151 =  n3149 & ~n3150;
assign n3152 =  n0338 & ~n0459;
assign n3153 =  n3151 & ~n3152;
assign n3154 =  n0339 & ~n0459;
assign n3155 =  n3153 & ~n3154;
assign n3156 =  n0453 & ~n0458;
assign n3157 =  n3155 & ~n3156;
assign n3158 =  n0457 & ~n0458;
assign n3159 =  n3157 & ~n3158;
assign n3160 =  n0336 & ~n0458;
assign n3161 =  n3159 & ~n3160;
assign n3162 =  n0337 & ~n0458;
assign n3163 =  n3161 & ~n3162;
assign n3164 =  n0338 & ~n0458;
assign n3165 =  n3163 & ~n3164;
assign n3166 =  n0339 & ~n0458;
assign n3167 =  n3165 & ~n3166;
assign n3168 =  n0455 &  n0456;
assign n3169 =  n0454 &  n3168;
assign n3170 = ~n0457 &  n3169;
assign n3171 =  n3167 & ~n3170;
assign n3172 =  n0396 & ~n0456;
assign n3173 =  n3171 & ~n3172;
assign n3174 =  n0379 & ~n0456;
assign n3175 =  n3173 & ~n3174;
assign n3176 =  n0397 & ~n0456;
assign n3177 =  n3175 & ~n3176;
assign n3178 =  n0380 & ~n0456;
assign n3179 =  n3177 & ~n3178;
assign n3180 =  n0381 & ~n0456;
assign n3181 =  n3179 & ~n3180;
assign n3182 =  n0398 & ~n0456;
assign n3183 =  n3181 & ~n3182;
assign n3184 =  n0399 & ~n0456;
assign n3185 =  n3183 & ~n3184;
assign n3186 =  n0076 & ~n0456;
assign n3187 =  n3185 & ~n3186;
assign n3188 =  n0073 & ~n0456;
assign n3189 =  n3187 & ~n3188;
assign n3190 =  n0069 & ~n0456;
assign n3191 =  n3189 & ~n3190;
assign n3192 =  n0068 & ~n0456;
assign n3193 =  n3191 & ~n3192;
assign n3194 =  n0054 & ~n0456;
assign n3195 =  n3193 & ~n3194;
assign n3196 =  n0053 & ~n0456;
assign n3197 =  n3195 & ~n3196;
assign n3198 =  n0052 & ~n0456;
assign n3199 =  n3197 & ~n3198;
assign n3200 =  n0382 & ~n0456;
assign n3201 =  n3199 & ~n3200;
assign n3202 =  n0391 & ~n0455;
assign n3203 =  n3201 & ~n3202;
assign n3204 =  n0374 & ~n0455;
assign n3205 =  n3203 & ~n3204;
assign n3206 =  n0392 & ~n0455;
assign n3207 =  n3205 & ~n3206;
assign n3208 =  n0375 & ~n0455;
assign n3209 =  n3207 & ~n3208;
assign n3210 =  n0393 & ~n0455;
assign n3211 =  n3209 & ~n3210;
assign n3212 =  n0394 & ~n0455;
assign n3213 =  n3211 & ~n3212;
assign n3214 =  n0376 & ~n0455;
assign n3215 =  n3213 & ~n3214;
assign n3216 =  n0075 & ~n0455;
assign n3217 =  n3215 & ~n3216;
assign n3218 =  n0072 & ~n0455;
assign n3219 =  n3217 & ~n3218;
assign n3220 =  n0066 & ~n0455;
assign n3221 =  n3219 & ~n3220;
assign n3222 =  n0065 & ~n0455;
assign n3223 =  n3221 & ~n3222;
assign n3224 =  n0041 & ~n0455;
assign n3225 =  n3223 & ~n3224;
assign n3226 =  n0040 & ~n0455;
assign n3227 =  n3225 & ~n3226;
assign n3228 =  n0377 & ~n0455;
assign n3229 =  n3227 & ~n3228;
assign n3230 =  n0039 & ~n0455;
assign n3231 =  n3229 & ~n3230;
assign n3232 =  n0386 & ~n0454;
assign n3233 =  n3231 & ~n3232;
assign n3234 =  n0387 & ~n0454;
assign n3235 =  n3233 & ~n3234;
assign n3236 =  n0369 & ~n0454;
assign n3237 =  n3235 & ~n3236;
assign n3238 =  n0388 & ~n0454;
assign n3239 =  n3237 & ~n3238;
assign n3240 =  n0389 & ~n0454;
assign n3241 =  n3239 & ~n3240;
assign n3242 =  n0370 & ~n0454;
assign n3243 =  n3241 & ~n3242;
assign n3244 =  n0371 & ~n0454;
assign n3245 =  n3243 & ~n3244;
assign n3246 =  n0372 & ~n0454;
assign n3247 =  n3245 & ~n3246;
assign n3248 =  n0074 & ~n0454;
assign n3249 =  n3247 & ~n3248;
assign n3250 =  n0071 & ~n0454;
assign n3251 =  n3249 & ~n3250;
assign n3252 =  n0063 & ~n0454;
assign n3253 =  n3251 & ~n3252;
assign n3254 =  n0062 & ~n0454;
assign n3255 =  n3253 & ~n3254;
assign n3256 =  n0028 & ~n0454;
assign n3257 =  n3255 & ~n3256;
assign n3258 =  n0027 & ~n0454;
assign n3259 =  n3257 & ~n3258;
assign n3260 =  n0026 & ~n0454;
assign n3261 =  n3259 & ~n3260;
assign n3262 = ~n0453 &  n2663;
assign n3263 =  n3261 & ~n3262;
assign n3264 =  n0417 & ~n0452;
assign n3265 =  n3263 & ~n3264;
assign n3266 =  n0336 & ~n0452;
assign n3267 =  n3265 & ~n3266;
assign n3268 =  n0337 & ~n0452;
assign n3269 =  n3267 & ~n3268;
assign n3270 =  n0338 & ~n0452;
assign n3271 =  n3269 & ~n3270;
assign n3272 =  n0339 & ~n0452;
assign n3273 =  n3271 & ~n3272;
assign n3274 =  n0422 & ~n0451;
assign n3275 =  n3273 & ~n3274;
assign n3276 =  n0450 & ~n0451;
assign n3277 =  n3275 & ~n3276;
assign n3278 =  n0336 & ~n0451;
assign n3279 =  n3277 & ~n3278;
assign n3280 =  n0337 & ~n0451;
assign n3281 =  n3279 & ~n3280;
assign n3282 =  n0338 & ~n0451;
assign n3283 =  n3281 & ~n3282;
assign n3284 =  n0339 & ~n0451;
assign n3285 =  n3283 & ~n3284;
assign n3286 =  n0448 &  n0449;
assign n3287 =  n0447 &  n3286;
assign n3288 = ~n0450 &  n3287;
assign n3289 =  n3285 & ~n3288;
assign n3290 =  n0412 & ~n0449;
assign n3291 =  n3289 & ~n3290;
assign n3292 =  n0435 & ~n0449;
assign n3293 =  n3291 & ~n3292;
assign n3294 =  n0436 & ~n0449;
assign n3295 =  n3293 & ~n3294;
assign n3296 =  n0413 & ~n0449;
assign n3297 =  n3295 & ~n3296;
assign n3298 =  n0414 & ~n0449;
assign n3299 =  n3297 & ~n3298;
assign n3300 =  n0437 & ~n0449;
assign n3301 =  n3299 & ~n3300;
assign n3302 =  n0438 & ~n0449;
assign n3303 =  n3301 & ~n3302;
assign n3304 =  n0415 & ~n0449;
assign n3305 =  n3303 & ~n3304;
assign n3306 =  n0076 & ~n0449;
assign n3307 =  n3305 & ~n3306;
assign n3308 =  n0073 & ~n0449;
assign n3309 =  n3307 & ~n3308;
assign n3310 =  n0068 & ~n0449;
assign n3311 =  n3309 & ~n3310;
assign n3312 =  n0054 & ~n0449;
assign n3313 =  n3311 & ~n3312;
assign n3314 =  n0053 & ~n0449;
assign n3315 =  n3313 & ~n3314;
assign n3316 =  n0052 & ~n0449;
assign n3317 =  n3315 & ~n3316;
assign n3318 =  n0051 & ~n0449;
assign n3319 =  n3317 & ~n3318;
assign n3320 =  n0430 & ~n0448;
assign n3321 =  n3319 & ~n3320;
assign n3322 =  n0431 & ~n0448;
assign n3323 =  n3321 & ~n3322;
assign n3324 =  n0432 & ~n0448;
assign n3325 =  n3323 & ~n3324;
assign n3326 =  n0407 & ~n0448;
assign n3327 =  n3325 & ~n3326;
assign n3328 =  n0433 & ~n0448;
assign n3329 =  n3327 & ~n3328;
assign n3330 =  n0408 & ~n0448;
assign n3331 =  n3329 & ~n3330;
assign n3332 =  n0409 & ~n0448;
assign n3333 =  n3331 & ~n3332;
assign n3334 =  n0410 & ~n0448;
assign n3335 =  n3333 & ~n3334;
assign n3336 =  n0075 & ~n0448;
assign n3337 =  n3335 & ~n3336;
assign n3338 =  n0072 & ~n0448;
assign n3339 =  n3337 & ~n3338;
assign n3340 =  n0065 & ~n0448;
assign n3341 =  n3339 & ~n3340;
assign n3342 =  n0041 & ~n0448;
assign n3343 =  n3341 & ~n3342;
assign n3344 =  n0040 & ~n0448;
assign n3345 =  n3343 & ~n3344;
assign n3346 =  n0039 & ~n0448;
assign n3347 =  n3345 & ~n3346;
assign n3348 =  n0038 & ~n0448;
assign n3349 =  n3347 & ~n3348;
assign n3350 =  n0402 & ~n0447;
assign n3351 =  n3349 & ~n3350;
assign n3352 =  n0425 & ~n0447;
assign n3353 =  n3351 & ~n3352;
assign n3354 =  n0426 & ~n0447;
assign n3355 =  n3353 & ~n3354;
assign n3356 =  n0427 & ~n0447;
assign n3357 =  n3355 & ~n3356;
assign n3358 =  n0403 & ~n0447;
assign n3359 =  n3357 & ~n3358;
assign n3360 =  n0404 & ~n0447;
assign n3361 =  n3359 & ~n3360;
assign n3362 =  n0405 & ~n0447;
assign n3363 =  n3361 & ~n3362;
assign n3364 =  n0074 & ~n0447;
assign n3365 =  n3363 & ~n3364;
assign n3366 =  n0071 & ~n0447;
assign n3367 =  n3365 & ~n3366;
assign n3368 =  n0062 & ~n0447;
assign n3369 =  n3367 & ~n3368;
assign n3370 =  n0428 & ~n0447;
assign n3371 =  n3369 & ~n3370;
assign n3372 =  n0028 & ~n0447;
assign n3373 =  n3371 & ~n3372;
assign n3374 =  n0027 & ~n0447;
assign n3375 =  n3373 & ~n3374;
assign n3376 =  n0026 & ~n0447;
assign n3377 =  n3375 & ~n3376;
assign n3378 =  n0025 & ~n0447;
assign n3379 =  n3377 & ~n3378;
assign n3380 =  n0384 & ~n0446;
assign n3381 =  n3379 & ~n3380;
assign n3382 =  n0445 & ~n0446;
assign n3383 =  n3381 & ~n3382;
assign n3384 =  n0336 & ~n0446;
assign n3385 =  n3383 & ~n3384;
assign n3386 =  n0337 & ~n0446;
assign n3387 =  n3385 & ~n3386;
assign n3388 =  n0338 & ~n0446;
assign n3389 =  n3387 & ~n3388;
assign n3390 =  n0339 & ~n0446;
assign n3391 =  n3389 & ~n3390;
assign n3392 =  n0443 &  n0444;
assign n3393 =  n0442 &  n3392;
assign n3394 = ~n0445 &  n3393;
assign n3395 =  n3391 & ~n3394;
assign n3396 =  n0360 & ~n0444;
assign n3397 =  n3395 & ~n3396;
assign n3398 =  n0412 & ~n0444;
assign n3399 =  n3397 & ~n3398;
assign n3400 =  n0361 & ~n0444;
assign n3401 =  n3399 & ~n3400;
assign n3402 =  n0364 & ~n0444;
assign n3403 =  n3401 & ~n3402;
assign n3404 =  n0413 & ~n0444;
assign n3405 =  n3403 & ~n3404;
assign n3406 =  n0366 & ~n0444;
assign n3407 =  n3405 & ~n3406;
assign n3408 =  n0414 & ~n0444;
assign n3409 =  n3407 & ~n3408;
assign n3410 =  n0415 & ~n0444;
assign n3411 =  n3409 & ~n3410;
assign n3412 =  n0073 & ~n0444;
assign n3413 =  n3411 & ~n3412;
assign n3414 =  n0070 & ~n0444;
assign n3415 =  n3413 & ~n3414;
assign n3416 =  n0069 & ~n0444;
assign n3417 =  n3415 & ~n3416;
assign n3418 =  n0068 & ~n0444;
assign n3419 =  n3417 & ~n3418;
assign n3420 =  n0055 & ~n0444;
assign n3421 =  n3419 & ~n3420;
assign n3422 =  n0053 & ~n0444;
assign n3423 =  n3421 & ~n3422;
assign n3424 =  n0052 & ~n0444;
assign n3425 =  n3423 & ~n3424;
assign n3426 =  n0350 & ~n0443;
assign n3427 =  n3425 & ~n3426;
assign n3428 =  n0351 & ~n0443;
assign n3429 =  n3427 & ~n3428;
assign n3430 =  n0353 & ~n0443;
assign n3431 =  n3429 & ~n3430;
assign n3432 =  n0355 & ~n0443;
assign n3433 =  n3431 & ~n3432;
assign n3434 =  n0407 & ~n0443;
assign n3435 =  n3433 & ~n3434;
assign n3436 =  n0408 & ~n0443;
assign n3437 =  n3435 & ~n3436;
assign n3438 =  n0409 & ~n0443;
assign n3439 =  n3437 & ~n3438;
assign n3440 =  n0410 & ~n0443;
assign n3441 =  n3439 & ~n3440;
assign n3442 =  n0072 & ~n0443;
assign n3443 =  n3441 & ~n3442;
assign n3444 =  n0067 & ~n0443;
assign n3445 =  n3443 & ~n3444;
assign n3446 =  n0066 & ~n0443;
assign n3447 =  n3445 & ~n3446;
assign n3448 =  n0065 & ~n0443;
assign n3449 =  n3447 & ~n3448;
assign n3450 =  n0042 & ~n0443;
assign n3451 =  n3449 & ~n3450;
assign n3452 =  n0040 & ~n0443;
assign n3453 =  n3451 & ~n3452;
assign n3454 =  n0039 & ~n0443;
assign n3455 =  n3453 & ~n3454;
assign n3456 =  n0342 & ~n0442;
assign n3457 =  n3455 & ~n3456;
assign n3458 =  n0343 & ~n0442;
assign n3459 =  n3457 & ~n3458;
assign n3460 =  n0344 & ~n0442;
assign n3461 =  n3459 & ~n3460;
assign n3462 =  n0402 & ~n0442;
assign n3463 =  n3461 & ~n3462;
assign n3464 =  n0403 & ~n0442;
assign n3465 =  n3463 & ~n3464;
assign n3466 =  n0404 & ~n0442;
assign n3467 =  n3465 & ~n3466;
assign n3468 =  n0347 & ~n0442;
assign n3469 =  n3467 & ~n3468;
assign n3470 =  n0405 & ~n0442;
assign n3471 =  n3469 & ~n3470;
assign n3472 =  n0071 & ~n0442;
assign n3473 =  n3471 & ~n3472;
assign n3474 =  n0064 & ~n0442;
assign n3475 =  n3473 & ~n3474;
assign n3476 =  n0063 & ~n0442;
assign n3477 =  n3475 & ~n3476;
assign n3478 =  n0062 & ~n0442;
assign n3479 =  n3477 & ~n3478;
assign n3480 =  n0029 & ~n0442;
assign n3481 =  n3479 & ~n3480;
assign n3482 =  n0027 & ~n0442;
assign n3483 =  n3481 & ~n3482;
assign n3484 =  n0026 & ~n0442;
assign n3485 =  n3483 & ~n3484;
assign n3486 =  n0424 & ~n0441;
assign n3487 =  n3485 & ~n3486;
assign n3488 =  n0440 & ~n0441;
assign n3489 =  n3487 & ~n3488;
assign n3490 =  n0336 & ~n0441;
assign n3491 =  n3489 & ~n3490;
assign n3492 =  n0337 & ~n0441;
assign n3493 =  n3491 & ~n3492;
assign n3494 =  n0338 & ~n0441;
assign n3495 =  n3493 & ~n3494;
assign n3496 =  n0339 & ~n0441;
assign n3497 =  n3495 & ~n3496;
assign n3498 =  n0434 &  n0439;
assign n3499 =  n0429 &  n3498;
assign n3500 = ~n0440 &  n3499;
assign n3501 =  n3497 & ~n3500;
assign n3502 =  n0379 & ~n0439;
assign n3503 =  n3501 & ~n3502;
assign n3504 =  n0435 & ~n0439;
assign n3505 =  n3503 & ~n3504;
assign n3506 =  n0436 & ~n0439;
assign n3507 =  n3505 & ~n3506;
assign n3508 =  n0380 & ~n0439;
assign n3509 =  n3507 & ~n3508;
assign n3510 =  n0437 & ~n0439;
assign n3511 =  n3509 & ~n3510;
assign n3512 =  n0381 & ~n0439;
assign n3513 =  n3511 & ~n3512;
assign n3514 =  n0438 & ~n0439;
assign n3515 =  n3513 & ~n3514;
assign n3516 =  n0073 & ~n0439;
assign n3517 =  n3515 & ~n3516;
assign n3518 =  n0068 & ~n0439;
assign n3519 =  n3517 & ~n3518;
assign n3520 =  n0055 & ~n0439;
assign n3521 =  n3519 & ~n3520;
assign n3522 =  n0054 & ~n0439;
assign n3523 =  n3521 & ~n3522;
assign n3524 =  n0053 & ~n0439;
assign n3525 =  n3523 & ~n3524;
assign n3526 =  n0052 & ~n0439;
assign n3527 =  n3525 & ~n3526;
assign n3528 =  n0051 & ~n0439;
assign n3529 =  n3527 & ~n3528;
assign n3530 =  n0382 & ~n0439;
assign n3531 =  n3529 & ~n3530;
assign n3532 =  n0010 &  n0061;
assign n3533 = ~n0438 &  n3532;
assign n3534 =  n3531 & ~n3533;
assign n3535 = ~n0009 &  n0057;
assign n3536 = ~n0437 &  n3535;
assign n3537 =  n3534 & ~n3536;
assign n3538 =  n0009 &  n0059;
assign n3539 = ~n0436 &  n3538;
assign n3540 =  n3537 & ~n3539;
assign n3541 = ~n0010 &  n0058;
assign n3542 = ~n0435 &  n3541;
assign n3543 =  n3540 & ~n3542;
assign n3544 =  n0430 & ~n0434;
assign n3545 =  n3543 & ~n3544;
assign n3546 =  n0431 & ~n0434;
assign n3547 =  n3545 & ~n3546;
assign n3548 =  n0432 & ~n0434;
assign n3549 =  n3547 & ~n3548;
assign n3550 =  n0374 & ~n0434;
assign n3551 =  n3549 & ~n3550;
assign n3552 =  n0375 & ~n0434;
assign n3553 =  n3551 & ~n3552;
assign n3554 =  n0433 & ~n0434;
assign n3555 =  n3553 & ~n3554;
assign n3556 =  n0376 & ~n0434;
assign n3557 =  n3555 & ~n3556;
assign n3558 =  n0072 & ~n0434;
assign n3559 =  n3557 & ~n3558;
assign n3560 =  n0065 & ~n0434;
assign n3561 =  n3559 & ~n3560;
assign n3562 =  n0042 & ~n0434;
assign n3563 =  n3561 & ~n3562;
assign n3564 =  n0041 & ~n0434;
assign n3565 =  n3563 & ~n3564;
assign n3566 =  n0040 & ~n0434;
assign n3567 =  n3565 & ~n3566;
assign n3568 =  n0377 & ~n0434;
assign n3569 =  n3567 & ~n3568;
assign n3570 =  n0039 & ~n0434;
assign n3571 =  n3569 & ~n3570;
assign n3572 =  n0038 & ~n0434;
assign n3573 =  n3571 & ~n3572;
assign n3574 = ~n0009 &  n0044;
assign n3575 = ~n0433 &  n3574;
assign n3576 =  n3573 & ~n3575;
assign n3577 =  n0009 &  n0046;
assign n3578 = ~n0432 &  n3577;
assign n3579 =  n3576 & ~n3578;
assign n3580 =  n0010 &  n0048;
assign n3581 = ~n0431 &  n3580;
assign n3582 =  n3579 & ~n3581;
assign n3583 = ~n0010 &  n0045;
assign n3584 = ~n0430 &  n3583;
assign n3585 =  n3582 & ~n3584;
assign n3586 =  n0425 & ~n0429;
assign n3587 =  n3585 & ~n3586;
assign n3588 =  n0426 & ~n0429;
assign n3589 =  n3587 & ~n3588;
assign n3590 =  n0369 & ~n0429;
assign n3591 =  n3589 & ~n3590;
assign n3592 =  n0427 & ~n0429;
assign n3593 =  n3591 & ~n3592;
assign n3594 =  n0370 & ~n0429;
assign n3595 =  n3593 & ~n3594;
assign n3596 =  n0371 & ~n0429;
assign n3597 =  n3595 & ~n3596;
assign n3598 =  n0372 & ~n0429;
assign n3599 =  n3597 & ~n3598;
assign n3600 =  n0071 & ~n0429;
assign n3601 =  n3599 & ~n3600;
assign n3602 =  n0062 & ~n0429;
assign n3603 =  n3601 & ~n3602;
assign n3604 =  n0428 & ~n0429;
assign n3605 =  n3603 & ~n3604;
assign n3606 =  n0029 & ~n0429;
assign n3607 =  n3605 & ~n3606;
assign n3608 =  n0028 & ~n0429;
assign n3609 =  n3607 & ~n3608;
assign n3610 =  n0027 & ~n0429;
assign n3611 =  n3609 & ~n3610;
assign n3612 =  n0026 & ~n0429;
assign n3613 =  n3611 & ~n3612;
assign n3614 =  n0025 & ~n0429;
assign n3615 =  n3613 & ~n3614;
assign n3616 =  n0009 &  n0033;
assign n3617 = ~n0428 &  n3616;
assign n3618 =  n3615 & ~n3617;
assign n3619 = ~n0009 &  n0031;
assign n3620 = ~n0427 &  n3619;
assign n3621 =  n3618 & ~n3620;
assign n3622 =  n0010 &  n0035;
assign n3623 = ~n0426 &  n3622;
assign n3624 =  n3621 & ~n3623;
assign n3625 = ~n0010 &  n0032;
assign n3626 = ~n0425 &  n3625;
assign n3627 =  n3624 & ~n3626;
assign n3628 =  n0418 &  n0423;
assign n3629 =  n0385 &  n3628;
assign n3630 = ~n0424 &  n3629;
assign n3631 =  n3627 & ~n3630;
assign n3632 =  n0422 & ~n0423;
assign n3633 =  n3631 & ~n3632;
assign n3634 =  n0336 & ~n0423;
assign n3635 =  n3633 & ~n3634;
assign n3636 =  n0337 & ~n0423;
assign n3637 =  n3635 & ~n3636;
assign n3638 =  n0338 & ~n0423;
assign n3639 =  n3637 & ~n3638;
assign n3640 =  n0339 & ~n0423;
assign n3641 =  n3639 & ~n3640;
assign n3642 =  n0420 &  n0421;
assign n3643 =  n0419 &  n3642;
assign n3644 = ~n0422 &  n3643;
assign n3645 =  n3641 & ~n3644;
assign n3646 =  n0359 & ~n0421;
assign n3647 =  n3645 & ~n3646;
assign n3648 =  n0326 & ~n0421;
assign n3649 =  n3647 & ~n3648;
assign n3650 =  n0362 & ~n0421;
assign n3651 =  n3649 & ~n3650;
assign n3652 =  n0363 & ~n0421;
assign n3653 =  n3651 & ~n3652;
assign n3654 =  n0327 & ~n0421;
assign n3655 =  n3653 & ~n3654;
assign n3656 =  n0329 & ~n0421;
assign n3657 =  n3655 & ~n3656;
assign n3658 =  n0365 & ~n0421;
assign n3659 =  n3657 & ~n3658;
assign n3660 =  n0333 & ~n0421;
assign n3661 =  n3659 & ~n3660;
assign n3662 =  n0079 & ~n0421;
assign n3663 =  n3661 & ~n3662;
assign n3664 =  n0069 & ~n0421;
assign n3665 =  n3663 & ~n3664;
assign n3666 =  n0068 & ~n0421;
assign n3667 =  n3665 & ~n3666;
assign n3668 =  n0055 & ~n0421;
assign n3669 =  n3667 & ~n3668;
assign n3670 =  n0054 & ~n0421;
assign n3671 =  n3669 & ~n3670;
assign n3672 =  n0052 & ~n0421;
assign n3673 =  n3671 & ~n3672;
assign n3674 =  n0050 & ~n0421;
assign n3675 =  n3673 & ~n3674;
assign n3676 =  n0317 & ~n0420;
assign n3677 =  n3675 & ~n3676;
assign n3678 =  n0352 & ~n0420;
assign n3679 =  n3677 & ~n3678;
assign n3680 =  n0354 & ~n0420;
assign n3681 =  n3679 & ~n3680;
assign n3682 =  n0318 & ~n0420;
assign n3683 =  n3681 & ~n3682;
assign n3684 =  n0356 & ~n0420;
assign n3685 =  n3683 & ~n3684;
assign n3686 =  n0321 & ~n0420;
assign n3687 =  n3685 & ~n3686;
assign n3688 =  n0357 & ~n0420;
assign n3689 =  n3687 & ~n3688;
assign n3690 =  n0323 & ~n0420;
assign n3691 =  n3689 & ~n3690;
assign n3692 =  n0078 & ~n0420;
assign n3693 =  n3691 & ~n3692;
assign n3694 =  n0066 & ~n0420;
assign n3695 =  n3693 & ~n3694;
assign n3696 =  n0065 & ~n0420;
assign n3697 =  n3695 & ~n3696;
assign n3698 =  n0042 & ~n0420;
assign n3699 =  n3697 & ~n3698;
assign n3700 =  n0041 & ~n0420;
assign n3701 =  n3699 & ~n3700;
assign n3702 =  n0039 & ~n0420;
assign n3703 =  n3701 & ~n3702;
assign n3704 =  n0037 & ~n0420;
assign n3705 =  n3703 & ~n3704;
assign n3706 =  n0341 & ~n0419;
assign n3707 =  n3705 & ~n3706;
assign n3708 =  n0345 & ~n0419;
assign n3709 =  n3707 & ~n3708;
assign n3710 =  n0308 & ~n0419;
assign n3711 =  n3709 & ~n3710;
assign n3712 =  n0346 & ~n0419;
assign n3713 =  n3711 & ~n3712;
assign n3714 =  n0311 & ~n0419;
assign n3715 =  n3713 & ~n3714;
assign n3716 =  n0312 & ~n0419;
assign n3717 =  n3715 & ~n3716;
assign n3718 =  n0348 & ~n0419;
assign n3719 =  n3717 & ~n3718;
assign n3720 =  n0077 & ~n0419;
assign n3721 =  n3719 & ~n3720;
assign n3722 =  n0063 & ~n0419;
assign n3723 =  n3721 & ~n3722;
assign n3724 =  n0062 & ~n0419;
assign n3725 =  n3723 & ~n3724;
assign n3726 =  n0315 & ~n0419;
assign n3727 =  n3725 & ~n3726;
assign n3728 =  n0029 & ~n0419;
assign n3729 =  n3727 & ~n3728;
assign n3730 =  n0028 & ~n0419;
assign n3731 =  n3729 & ~n3730;
assign n3732 =  n0026 & ~n0419;
assign n3733 =  n3731 & ~n3732;
assign n3734 =  n0024 & ~n0419;
assign n3735 =  n3733 & ~n3734;
assign n3736 =  n0401 & ~n0418;
assign n3737 =  n3735 & ~n3736;
assign n3738 =  n0417 & ~n0418;
assign n3739 =  n3737 & ~n3738;
assign n3740 =  n0336 & ~n0418;
assign n3741 =  n3739 & ~n3740;
assign n3742 =  n0337 & ~n0418;
assign n3743 =  n3741 & ~n3742;
assign n3744 =  n0338 & ~n0418;
assign n3745 =  n3743 & ~n3744;
assign n3746 =  n0339 & ~n0418;
assign n3747 =  n3745 & ~n3746;
assign n3748 =  n0411 &  n0416;
assign n3749 =  n0406 &  n3748;
assign n3750 = ~n0417 &  n3749;
assign n3751 =  n3747 & ~n3750;
assign n3752 =  n0326 & ~n0416;
assign n3753 =  n3751 & ~n3752;
assign n3754 =  n0412 & ~n0416;
assign n3755 =  n3753 & ~n3754;
assign n3756 =  n0327 & ~n0416;
assign n3757 =  n3755 & ~n3756;
assign n3758 =  n0329 & ~n0416;
assign n3759 =  n3757 & ~n3758;
assign n3760 =  n0413 & ~n0416;
assign n3761 =  n3759 & ~n3760;
assign n3762 =  n0414 & ~n0416;
assign n3763 =  n3761 & ~n3762;
assign n3764 =  n0333 & ~n0416;
assign n3765 =  n3763 & ~n3764;
assign n3766 =  n0415 & ~n0416;
assign n3767 =  n3765 & ~n3766;
assign n3768 =  n0079 & ~n0416;
assign n3769 =  n3767 & ~n3768;
assign n3770 =  n0073 & ~n0416;
assign n3771 =  n3769 & ~n3770;
assign n3772 =  n0069 & ~n0416;
assign n3773 =  n3771 & ~n3772;
assign n3774 =  n0068 & ~n0416;
assign n3775 =  n3773 & ~n3774;
assign n3776 =  n0055 & ~n0416;
assign n3777 =  n3775 & ~n3776;
assign n3778 =  n0054 & ~n0416;
assign n3779 =  n3777 & ~n3778;
assign n3780 =  n0052 & ~n0416;
assign n3781 =  n3779 & ~n3780;
assign n3782 =  n0011 &  n0022;
assign n3783 = ~n0415 &  n3782;
assign n3784 =  n3781 & ~n3783;
assign n3785 =  n0012 &  n0060;
assign n3786 = ~n0414 &  n3785;
assign n3787 =  n3784 & ~n3786;
assign n3788 = ~n0011 &  n0019;
assign n3789 = ~n0413 &  n3788;
assign n3790 =  n3787 & ~n3789;
assign n3791 = ~n0012 &  n0056;
assign n3792 = ~n0412 &  n3791;
assign n3793 =  n3790 & ~n3792;
assign n3794 =  n0317 & ~n0411;
assign n3795 =  n3793 & ~n3794;
assign n3796 =  n0318 & ~n0411;
assign n3797 =  n3795 & ~n3796;
assign n3798 =  n0407 & ~n0411;
assign n3799 =  n3797 & ~n3798;
assign n3800 =  n0321 & ~n0411;
assign n3801 =  n3799 & ~n3800;
assign n3802 =  n0408 & ~n0411;
assign n3803 =  n3801 & ~n3802;
assign n3804 =  n0409 & ~n0411;
assign n3805 =  n3803 & ~n3804;
assign n3806 =  n0410 & ~n0411;
assign n3807 =  n3805 & ~n3806;
assign n3808 =  n0323 & ~n0411;
assign n3809 =  n3807 & ~n3808;
assign n3810 =  n0078 & ~n0411;
assign n3811 =  n3809 & ~n3810;
assign n3812 =  n0072 & ~n0411;
assign n3813 =  n3811 & ~n3812;
assign n3814 =  n0066 & ~n0411;
assign n3815 =  n3813 & ~n3814;
assign n3816 =  n0065 & ~n0411;
assign n3817 =  n3815 & ~n3816;
assign n3818 =  n0042 & ~n0411;
assign n3819 =  n3817 & ~n3818;
assign n3820 =  n0041 & ~n0411;
assign n3821 =  n3819 & ~n3820;
assign n3822 =  n0039 & ~n0411;
assign n3823 =  n3821 & ~n3822;
assign n3824 =  n0011 &  n0020;
assign n3825 = ~n0410 &  n3824;
assign n3826 =  n3823 & ~n3825;
assign n3827 =  n0012 &  n0047;
assign n3828 = ~n0409 &  n3827;
assign n3829 =  n3826 & ~n3828;
assign n3830 = ~n0012 &  n0043;
assign n3831 = ~n0408 &  n3830;
assign n3832 =  n3829 & ~n3831;
assign n3833 = ~n0011 &  n0018;
assign n3834 = ~n0407 &  n3833;
assign n3835 =  n3832 & ~n3834;
assign n3836 =  n0402 & ~n0406;
assign n3837 =  n3835 & ~n3836;
assign n3838 =  n0308 & ~n0406;
assign n3839 =  n3837 & ~n3838;
assign n3840 =  n0403 & ~n0406;
assign n3841 =  n3839 & ~n3840;
assign n3842 =  n0311 & ~n0406;
assign n3843 =  n3841 & ~n3842;
assign n3844 =  n0312 & ~n0406;
assign n3845 =  n3843 & ~n3844;
assign n3846 =  n0404 & ~n0406;
assign n3847 =  n3845 & ~n3846;
assign n3848 =  n0405 & ~n0406;
assign n3849 =  n3847 & ~n3848;
assign n3850 =  n0077 & ~n0406;
assign n3851 =  n3849 & ~n3850;
assign n3852 =  n0071 & ~n0406;
assign n3853 =  n3851 & ~n3852;
assign n3854 =  n0063 & ~n0406;
assign n3855 =  n3853 & ~n3854;
assign n3856 =  n0062 & ~n0406;
assign n3857 =  n3855 & ~n3856;
assign n3858 =  n0315 & ~n0406;
assign n3859 =  n3857 & ~n3858;
assign n3860 =  n0029 & ~n0406;
assign n3861 =  n3859 & ~n3860;
assign n3862 =  n0028 & ~n0406;
assign n3863 =  n3861 & ~n3862;
assign n3864 =  n0026 & ~n0406;
assign n3865 =  n3863 & ~n3864;
assign n3866 =  n0011 &  n0021;
assign n3867 = ~n0405 &  n3866;
assign n3868 =  n3865 & ~n3867;
assign n3869 = ~n0011 &  n0017;
assign n3870 = ~n0404 &  n3869;
assign n3871 =  n3868 & ~n3870;
assign n3872 =  n0012 &  n0034;
assign n3873 = ~n0403 &  n3872;
assign n3874 =  n3871 & ~n3873;
assign n3875 = ~n0012 &  n0030;
assign n3876 = ~n0402 &  n3875;
assign n3877 =  n3874 & ~n3876;
assign n3878 =  n0395 &  n0400;
assign n3879 =  n0390 &  n3878;
assign n3880 = ~n0401 &  n3879;
assign n3881 =  n3877 & ~n3880;
assign n3882 =  n0359 & ~n0400;
assign n3883 =  n3881 & ~n3882;
assign n3884 =  n0396 & ~n0400;
assign n3885 =  n3883 & ~n3884;
assign n3886 =  n0362 & ~n0400;
assign n3887 =  n3885 & ~n3886;
assign n3888 =  n0363 & ~n0400;
assign n3889 =  n3887 & ~n3888;
assign n3890 =  n0397 & ~n0400;
assign n3891 =  n3889 & ~n3890;
assign n3892 =  n0365 & ~n0400;
assign n3893 =  n3891 & ~n3892;
assign n3894 =  n0398 & ~n0400;
assign n3895 =  n3893 & ~n3894;
assign n3896 =  n0399 & ~n0400;
assign n3897 =  n3895 & ~n3896;
assign n3898 =  n0070 & ~n0400;
assign n3899 =  n3897 & ~n3898;
assign n3900 =  n0069 & ~n0400;
assign n3901 =  n3899 & ~n3900;
assign n3902 =  n0068 & ~n0400;
assign n3903 =  n3901 & ~n3902;
assign n3904 =  n0055 & ~n0400;
assign n3905 =  n3903 & ~n3904;
assign n3906 =  n0053 & ~n0400;
assign n3907 =  n3905 & ~n3906;
assign n3908 =  n0052 & ~n0400;
assign n3909 =  n3907 & ~n3908;
assign n3910 =  n0050 & ~n0400;
assign n3911 =  n3909 & ~n3910;
assign n3912 =  n0012 &  n0061;
assign n3913 = ~n0399 &  n3912;
assign n3914 =  n3911 & ~n3913;
assign n3915 =  n0011 &  n0059;
assign n3916 = ~n0398 &  n3915;
assign n3917 =  n3914 & ~n3916;
assign n3918 = ~n0011 &  n0057;
assign n3919 = ~n0397 &  n3918;
assign n3920 =  n3917 & ~n3919;
assign n3921 = ~n0012 &  n0058;
assign n3922 = ~n0396 &  n3921;
assign n3923 =  n3920 & ~n3922;
assign n3924 =  n0391 & ~n0395;
assign n3925 =  n3923 & ~n3924;
assign n3926 =  n0352 & ~n0395;
assign n3927 =  n3925 & ~n3926;
assign n3928 =  n0354 & ~n0395;
assign n3929 =  n3927 & ~n3928;
assign n3930 =  n0356 & ~n0395;
assign n3931 =  n3929 & ~n3930;
assign n3932 =  n0392 & ~n0395;
assign n3933 =  n3931 & ~n3932;
assign n3934 =  n0357 & ~n0395;
assign n3935 =  n3933 & ~n3934;
assign n3936 =  n0393 & ~n0395;
assign n3937 =  n3935 & ~n3936;
assign n3938 =  n0394 & ~n0395;
assign n3939 =  n3937 & ~n3938;
assign n3940 =  n0067 & ~n0395;
assign n3941 =  n3939 & ~n3940;
assign n3942 =  n0066 & ~n0395;
assign n3943 =  n3941 & ~n3942;
assign n3944 =  n0065 & ~n0395;
assign n3945 =  n3943 & ~n3944;
assign n3946 =  n0042 & ~n0395;
assign n3947 =  n3945 & ~n3946;
assign n3948 =  n0040 & ~n0395;
assign n3949 =  n3947 & ~n3948;
assign n3950 =  n0039 & ~n0395;
assign n3951 =  n3949 & ~n3950;
assign n3952 =  n0037 & ~n0395;
assign n3953 =  n3951 & ~n3952;
assign n3954 =  n0012 &  n0048;
assign n3955 = ~n0394 &  n3954;
assign n3956 =  n3953 & ~n3955;
assign n3957 = ~n0011 &  n0044;
assign n3958 = ~n0393 &  n3957;
assign n3959 =  n3956 & ~n3958;
assign n3960 =  n0011 &  n0046;
assign n3961 = ~n0392 &  n3960;
assign n3962 =  n3959 & ~n3961;
assign n3963 = ~n0012 &  n0045;
assign n3964 = ~n0391 &  n3963;
assign n3965 =  n3962 & ~n3964;
assign n3966 =  n0341 & ~n0390;
assign n3967 =  n3965 & ~n3966;
assign n3968 =  n0386 & ~n0390;
assign n3969 =  n3967 & ~n3968;
assign n3970 =  n0387 & ~n0390;
assign n3971 =  n3969 & ~n3970;
assign n3972 =  n0345 & ~n0390;
assign n3973 =  n3971 & ~n3972;
assign n3974 =  n0346 & ~n0390;
assign n3975 =  n3973 & ~n3974;
assign n3976 =  n0388 & ~n0390;
assign n3977 =  n3975 & ~n3976;
assign n3978 =  n0389 & ~n0390;
assign n3979 =  n3977 & ~n3978;
assign n3980 =  n0348 & ~n0390;
assign n3981 =  n3979 & ~n3980;
assign n3982 =  n0064 & ~n0390;
assign n3983 =  n3981 & ~n3982;
assign n3984 =  n0063 & ~n0390;
assign n3985 =  n3983 & ~n3984;
assign n3986 =  n0062 & ~n0390;
assign n3987 =  n3985 & ~n3986;
assign n3988 =  n0029 & ~n0390;
assign n3989 =  n3987 & ~n3988;
assign n3990 =  n0027 & ~n0390;
assign n3991 =  n3989 & ~n3990;
assign n3992 =  n0026 & ~n0390;
assign n3993 =  n3991 & ~n3992;
assign n3994 =  n0024 & ~n0390;
assign n3995 =  n3993 & ~n3994;
assign n3996 = ~n0011 &  n0031;
assign n3997 = ~n0389 &  n3996;
assign n3998 =  n3995 & ~n3997;
assign n3999 =  n0011 &  n0033;
assign n4000 = ~n0388 &  n3999;
assign n4001 =  n3998 & ~n4000;
assign n4002 =  n0012 &  n0035;
assign n4003 = ~n0387 &  n4002;
assign n4004 =  n4001 & ~n4003;
assign n4005 = ~n0012 &  n0032;
assign n4006 = ~n0386 &  n4005;
assign n4007 =  n4004 & ~n4006;
assign n4008 =  n0368 & ~n0385;
assign n4009 =  n4007 & ~n4008;
assign n4010 =  n0384 & ~n0385;
assign n4011 =  n4009 & ~n4010;
assign n4012 =  n0336 & ~n0385;
assign n4013 =  n4011 & ~n4012;
assign n4014 =  n0337 & ~n0385;
assign n4015 =  n4013 & ~n4014;
assign n4016 =  n0338 & ~n0385;
assign n4017 =  n4015 & ~n4016;
assign n4018 =  n0339 & ~n0385;
assign n4019 =  n4017 & ~n4018;
assign n4020 =  n0378 &  n0383;
assign n4021 =  n0373 &  n4020;
assign n4022 = ~n0384 &  n4021;
assign n4023 =  n4019 & ~n4022;
assign n4024 =  n0326 & ~n0383;
assign n4025 =  n4023 & ~n4024;
assign n4026 =  n0379 & ~n0383;
assign n4027 =  n4025 & ~n4026;
assign n4028 =  n0327 & ~n0383;
assign n4029 =  n4027 & ~n4028;
assign n4030 =  n0329 & ~n0383;
assign n4031 =  n4029 & ~n4030;
assign n4032 =  n0380 & ~n0383;
assign n4033 =  n4031 & ~n4032;
assign n4034 =  n0381 & ~n0383;
assign n4035 =  n4033 & ~n4034;
assign n4036 =  n0333 & ~n0383;
assign n4037 =  n4035 & ~n4036;
assign n4038 =  n0079 & ~n0383;
assign n4039 =  n4037 & ~n4038;
assign n4040 =  n0073 & ~n0383;
assign n4041 =  n4039 & ~n4040;
assign n4042 =  n0070 & ~n0383;
assign n4043 =  n4041 & ~n4042;
assign n4044 =  n0069 & ~n0383;
assign n4045 =  n4043 & ~n4044;
assign n4046 =  n0068 & ~n0383;
assign n4047 =  n4045 & ~n4046;
assign n4048 =  n0055 & ~n0383;
assign n4049 =  n4047 & ~n4048;
assign n4050 =  n0052 & ~n0383;
assign n4051 =  n4049 & ~n4050;
assign n4052 =  n0382 & ~n0383;
assign n4053 =  n4051 & ~n4052;
assign n4054 = ~n0013 &  n0019;
assign n4055 = ~n0382 &  n4054;
assign n4056 =  n4053 & ~n4055;
assign n4057 =  n0013 &  n0022;
assign n4058 = ~n0381 &  n4057;
assign n4059 =  n4056 & ~n4058;
assign n4060 =  n0014 &  n0060;
assign n4061 = ~n0380 &  n4060;
assign n4062 =  n4059 & ~n4061;
assign n4063 = ~n0014 &  n0056;
assign n4064 = ~n0379 &  n4063;
assign n4065 =  n4062 & ~n4064;
assign n4066 =  n0317 & ~n0378;
assign n4067 =  n4065 & ~n4066;
assign n4068 =  n0318 & ~n0378;
assign n4069 =  n4067 & ~n4068;
assign n4070 =  n0374 & ~n0378;
assign n4071 =  n4069 & ~n4070;
assign n4072 =  n0321 & ~n0378;
assign n4073 =  n4071 & ~n4072;
assign n4074 =  n0375 & ~n0378;
assign n4075 =  n4073 & ~n4074;
assign n4076 =  n0376 & ~n0378;
assign n4077 =  n4075 & ~n4076;
assign n4078 =  n0323 & ~n0378;
assign n4079 =  n4077 & ~n4078;
assign n4080 =  n0078 & ~n0378;
assign n4081 =  n4079 & ~n4080;
assign n4082 =  n0072 & ~n0378;
assign n4083 =  n4081 & ~n4082;
assign n4084 =  n0067 & ~n0378;
assign n4085 =  n4083 & ~n4084;
assign n4086 =  n0066 & ~n0378;
assign n4087 =  n4085 & ~n4086;
assign n4088 =  n0065 & ~n0378;
assign n4089 =  n4087 & ~n4088;
assign n4090 =  n0042 & ~n0378;
assign n4091 =  n4089 & ~n4090;
assign n4092 =  n0377 & ~n0378;
assign n4093 =  n4091 & ~n4092;
assign n4094 =  n0039 & ~n0378;
assign n4095 =  n4093 & ~n4094;
assign n4096 =  n0013 &  n0020;
assign n4097 = ~n0377 &  n4096;
assign n4098 =  n4095 & ~n4097;
assign n4099 = ~n0013 &  n0018;
assign n4100 = ~n0376 &  n4099;
assign n4101 =  n4098 & ~n4100;
assign n4102 = ~n0014 &  n0043;
assign n4103 = ~n0375 &  n4102;
assign n4104 =  n4101 & ~n4103;
assign n4105 =  n0014 &  n0047;
assign n4106 = ~n0374 &  n4105;
assign n4107 =  n4104 & ~n4106;
assign n4108 =  n0308 & ~n0373;
assign n4109 =  n4107 & ~n4108;
assign n4110 =  n0369 & ~n0373;
assign n4111 =  n4109 & ~n4110;
assign n4112 =  n0311 & ~n0373;
assign n4113 =  n4111 & ~n4112;
assign n4114 =  n0312 & ~n0373;
assign n4115 =  n4113 & ~n4114;
assign n4116 =  n0370 & ~n0373;
assign n4117 =  n4115 & ~n4116;
assign n4118 =  n0371 & ~n0373;
assign n4119 =  n4117 & ~n4118;
assign n4120 =  n0372 & ~n0373;
assign n4121 =  n4119 & ~n4120;
assign n4122 =  n0077 & ~n0373;
assign n4123 =  n4121 & ~n4122;
assign n4124 =  n0071 & ~n0373;
assign n4125 =  n4123 & ~n4124;
assign n4126 =  n0064 & ~n0373;
assign n4127 =  n4125 & ~n4126;
assign n4128 =  n0063 & ~n0373;
assign n4129 =  n4127 & ~n4128;
assign n4130 =  n0062 & ~n0373;
assign n4131 =  n4129 & ~n4130;
assign n4132 =  n0315 & ~n0373;
assign n4133 =  n4131 & ~n4132;
assign n4134 =  n0029 & ~n0373;
assign n4135 =  n4133 & ~n4134;
assign n4136 =  n0026 & ~n0373;
assign n4137 =  n4135 & ~n4136;
assign n4138 =  n0014 &  n0034;
assign n4139 = ~n0372 &  n4138;
assign n4140 =  n4137 & ~n4139;
assign n4141 =  n0013 &  n0021;
assign n4142 = ~n0371 &  n4141;
assign n4143 =  n4140 & ~n4142;
assign n4144 = ~n0014 &  n0030;
assign n4145 = ~n0370 &  n4144;
assign n4146 =  n4143 & ~n4145;
assign n4147 = ~n0013 &  n0017;
assign n4148 = ~n0369 &  n4147;
assign n4149 =  n4146 & ~n4148;
assign n4150 =  n0358 &  n0367;
assign n4151 =  n0349 &  n4150;
assign n4152 = ~n0368 &  n4151;
assign n4153 =  n4149 & ~n4152;
assign n4154 =  n0359 & ~n0367;
assign n4155 =  n4153 & ~n4154;
assign n4156 =  n0360 & ~n0367;
assign n4157 =  n4155 & ~n4156;
assign n4158 =  n0361 & ~n0367;
assign n4159 =  n4157 & ~n4158;
assign n4160 =  n0362 & ~n0367;
assign n4161 =  n4159 & ~n4160;
assign n4162 =  n0363 & ~n0367;
assign n4163 =  n4161 & ~n4162;
assign n4164 =  n0364 & ~n0367;
assign n4165 =  n4163 & ~n4164;
assign n4166 =  n0365 & ~n0367;
assign n4167 =  n4165 & ~n4166;
assign n4168 =  n0366 & ~n0367;
assign n4169 =  n4167 & ~n4168;
assign n4170 =  n0069 & ~n0367;
assign n4171 =  n4169 & ~n4170;
assign n4172 =  n0068 & ~n0367;
assign n4173 =  n4171 & ~n4172;
assign n4174 =  n0055 & ~n0367;
assign n4175 =  n4173 & ~n4174;
assign n4176 =  n0054 & ~n0367;
assign n4177 =  n4175 & ~n4176;
assign n4178 =  n0053 & ~n0367;
assign n4179 =  n4177 & ~n4178;
assign n4180 =  n0052 & ~n0367;
assign n4181 =  n4179 & ~n4180;
assign n4182 =  n0050 & ~n0367;
assign n4183 =  n4181 & ~n4182;
assign n4184 =  n0014 &  n0061;
assign n4185 = ~n0366 &  n4184;
assign n4186 =  n4183 & ~n4185;
assign n4187 =  n0010 &  n0060;
assign n4188 = ~n0365 &  n4187;
assign n4189 =  n4186 & ~n4188;
assign n4190 = ~n0013 &  n0057;
assign n4191 = ~n0364 &  n4190;
assign n4192 =  n4189 & ~n4191;
assign n4193 =  n0009 &  n0022;
assign n4194 = ~n0363 &  n4193;
assign n4195 =  n4192 & ~n4194;
assign n4196 = ~n0009 &  n0019;
assign n4197 = ~n0362 &  n4196;
assign n4198 =  n4195 & ~n4197;
assign n4199 =  n0013 &  n0059;
assign n4200 = ~n0361 &  n4199;
assign n4201 =  n4198 & ~n4200;
assign n4202 = ~n0014 &  n0058;
assign n4203 = ~n0360 &  n4202;
assign n4204 =  n4201 & ~n4203;
assign n4205 = ~n0010 &  n0056;
assign n4206 = ~n0359 &  n4205;
assign n4207 =  n4204 & ~n4206;
assign n4208 =  n0350 & ~n0358;
assign n4209 =  n4207 & ~n4208;
assign n4210 =  n0351 & ~n0358;
assign n4211 =  n4209 & ~n4210;
assign n4212 =  n0352 & ~n0358;
assign n4213 =  n4211 & ~n4212;
assign n4214 =  n0353 & ~n0358;
assign n4215 =  n4213 & ~n4214;
assign n4216 =  n0354 & ~n0358;
assign n4217 =  n4215 & ~n4216;
assign n4218 =  n0355 & ~n0358;
assign n4219 =  n4217 & ~n4218;
assign n4220 =  n0356 & ~n0358;
assign n4221 =  n4219 & ~n4220;
assign n4222 =  n0357 & ~n0358;
assign n4223 =  n4221 & ~n4222;
assign n4224 =  n0066 & ~n0358;
assign n4225 =  n4223 & ~n4224;
assign n4226 =  n0065 & ~n0358;
assign n4227 =  n4225 & ~n4226;
assign n4228 =  n0042 & ~n0358;
assign n4229 =  n4227 & ~n4228;
assign n4230 =  n0041 & ~n0358;
assign n4231 =  n4229 & ~n4230;
assign n4232 =  n0040 & ~n0358;
assign n4233 =  n4231 & ~n4232;
assign n4234 =  n0039 & ~n0358;
assign n4235 =  n4233 & ~n4234;
assign n4236 =  n0037 & ~n0358;
assign n4237 =  n4235 & ~n4236;
assign n4238 =  n0009 &  n0020;
assign n4239 = ~n0357 &  n4238;
assign n4240 =  n4237 & ~n4239;
assign n4241 =  n0010 &  n0047;
assign n4242 = ~n0356 &  n4241;
assign n4243 =  n4240 & ~n4242;
assign n4244 = ~n0013 &  n0044;
assign n4245 = ~n0355 &  n4244;
assign n4246 =  n4243 & ~n4245;
assign n4247 = ~n0009 &  n0018;
assign n4248 = ~n0354 &  n4247;
assign n4249 =  n4246 & ~n4248;
assign n4250 =  n0013 &  n0046;
assign n4251 = ~n0353 &  n4250;
assign n4252 =  n4249 & ~n4251;
assign n4253 = ~n0010 &  n0043;
assign n4254 = ~n0352 &  n4253;
assign n4255 =  n4252 & ~n4254;
assign n4256 =  n0014 &  n0048;
assign n4257 = ~n0351 &  n4256;
assign n4258 =  n4255 & ~n4257;
assign n4259 = ~n0014 &  n0045;
assign n4260 = ~n0350 &  n4259;
assign n4261 =  n4258 & ~n4260;
assign n4262 =  n0341 & ~n0349;
assign n4263 =  n4261 & ~n4262;
assign n4264 =  n0342 & ~n0349;
assign n4265 =  n4263 & ~n4264;
assign n4266 =  n0343 & ~n0349;
assign n4267 =  n4265 & ~n4266;
assign n4268 =  n0344 & ~n0349;
assign n4269 =  n4267 & ~n4268;
assign n4270 =  n0345 & ~n0349;
assign n4271 =  n4269 & ~n4270;
assign n4272 =  n0346 & ~n0349;
assign n4273 =  n4271 & ~n4272;
assign n4274 =  n0347 & ~n0349;
assign n4275 =  n4273 & ~n4274;
assign n4276 =  n0348 & ~n0349;
assign n4277 =  n4275 & ~n4276;
assign n4278 =  n0063 & ~n0349;
assign n4279 =  n4277 & ~n4278;
assign n4280 =  n0062 & ~n0349;
assign n4281 =  n4279 & ~n4280;
assign n4282 =  n0029 & ~n0349;
assign n4283 =  n4281 & ~n4282;
assign n4284 =  n0028 & ~n0349;
assign n4285 =  n4283 & ~n4284;
assign n4286 =  n0027 & ~n0349;
assign n4287 =  n4285 & ~n4286;
assign n4288 =  n0026 & ~n0349;
assign n4289 =  n4287 & ~n4288;
assign n4290 =  n0024 & ~n0349;
assign n4291 =  n4289 & ~n4290;
assign n4292 =  n0009 &  n0021;
assign n4293 = ~n0348 &  n4292;
assign n4294 =  n4291 & ~n4293;
assign n4295 = ~n0013 &  n0031;
assign n4296 = ~n0347 &  n4295;
assign n4297 =  n4294 & ~n4296;
assign n4298 =  n0010 &  n0034;
assign n4299 = ~n0346 &  n4298;
assign n4300 =  n4297 & ~n4299;
assign n4301 = ~n0009 &  n0017;
assign n4302 = ~n0345 &  n4301;
assign n4303 =  n4300 & ~n4302;
assign n4304 =  n0014 &  n0035;
assign n4305 = ~n0344 &  n4304;
assign n4306 =  n4303 & ~n4305;
assign n4307 =  n0013 &  n0033;
assign n4308 = ~n0343 &  n4307;
assign n4309 =  n4306 & ~n4308;
assign n4310 = ~n0014 &  n0032;
assign n4311 = ~n0342 &  n4310;
assign n4312 =  n4309 & ~n4311;
assign n4313 = ~n0010 &  n0030;
assign n4314 = ~n0341 &  n4313;
assign n4315 =  n4312 & ~n4314;
assign n4316 =  n0335 & ~n0340;
assign n4317 =  n4315 & ~n4316;
assign n4318 =  n0336 & ~n0340;
assign n4319 =  n4317 & ~n4318;
assign n4320 =  n0337 & ~n0340;
assign n4321 =  n4319 & ~n4320;
assign n4322 =  n0338 & ~n0340;
assign n4323 =  n4321 & ~n4322;
assign n4324 =  n0339 & ~n0340;
assign n4325 =  n4323 & ~n4324;
assign n4326 = ~n0017 &  n0018;
assign n4327 = ~n0339 &  n4326;
assign n4328 =  n4325 & ~n4327;
assign n4329 = ~n0020 &  n0021;
assign n4330 = ~n0338 &  n4329;
assign n4331 =  n4328 & ~n4330;
assign n4332 = ~n0018 &  n0019;
assign n4333 = ~n0337 &  n4332;
assign n4334 =  n4331 & ~n4333;
assign n4335 =  n0020 & ~n0022;
assign n4336 = ~n0336 &  n4335;
assign n4337 =  n4334 & ~n4336;
assign n4338 =  n0325 &  n0334;
assign n4339 =  n0316 &  n4338;
assign n4340 = ~n0335 &  n4339;
assign n4341 =  n4337 & ~n4340;
assign n4342 =  n0326 & ~n0334;
assign n4343 =  n4341 & ~n4342;
assign n4344 =  n0327 & ~n0334;
assign n4345 =  n4343 & ~n4344;
assign n4346 =  n0328 & ~n0334;
assign n4347 =  n4345 & ~n4346;
assign n4348 =  n0329 & ~n0334;
assign n4349 =  n4347 & ~n4348;
assign n4350 =  n0330 & ~n0334;
assign n4351 =  n4349 & ~n4350;
assign n4352 =  n0331 & ~n0334;
assign n4353 =  n4351 & ~n4352;
assign n4354 =  n0332 & ~n0334;
assign n4355 =  n4353 & ~n4354;
assign n4356 =  n0333 & ~n0334;
assign n4357 =  n4355 & ~n4356;
assign n4358 =  n0082 & ~n0334;
assign n4359 =  n4357 & ~n4358;
assign n4360 =  n0079 & ~n0334;
assign n4361 =  n4359 & ~n4360;
assign n4362 =  n0073 & ~n0334;
assign n4363 =  n4361 & ~n4362;
assign n4364 =  n0069 & ~n0334;
assign n4365 =  n4363 & ~n4364;
assign n4366 =  n0055 & ~n0334;
assign n4367 =  n4365 & ~n4366;
assign n4368 =  n0054 & ~n0334;
assign n4369 =  n4367 & ~n4368;
assign n4370 =  n0049 & ~n0334;
assign n4371 =  n4369 & ~n4370;
assign n4372 =  n0016 &  n0061;
assign n4373 = ~n0333 &  n4372;
assign n4374 =  n4371 & ~n4373;
assign n4375 =  n0015 &  n0022;
assign n4376 = ~n0332 &  n4375;
assign n4377 =  n4374 & ~n4376;
assign n4378 =  n0016 &  n0060;
assign n4379 = ~n0331 &  n4378;
assign n4380 =  n4377 & ~n4379;
assign n4381 = ~n0016 &  n0056;
assign n4382 = ~n0330 &  n4381;
assign n4383 =  n4380 & ~n4382;
assign n4384 = ~n0016 &  n0058;
assign n4385 = ~n0329 &  n4384;
assign n4386 =  n4383 & ~n4385;
assign n4387 = ~n0015 &  n0019;
assign n4388 = ~n0328 &  n4387;
assign n4389 =  n4386 & ~n4388;
assign n4390 = ~n0015 &  n0057;
assign n4391 = ~n0327 &  n4390;
assign n4392 =  n4389 & ~n4391;
assign n4393 =  n0015 &  n0059;
assign n4394 = ~n0326 &  n4393;
assign n4395 =  n4392 & ~n4394;
assign n4396 =  n0317 & ~n0325;
assign n4397 =  n4395 & ~n4396;
assign n4398 =  n0318 & ~n0325;
assign n4399 =  n4397 & ~n4398;
assign n4400 =  n0319 & ~n0325;
assign n4401 =  n4399 & ~n4400;
assign n4402 =  n0320 & ~n0325;
assign n4403 =  n4401 & ~n4402;
assign n4404 =  n0321 & ~n0325;
assign n4405 =  n4403 & ~n4404;
assign n4406 =  n0322 & ~n0325;
assign n4407 =  n4405 & ~n4406;
assign n4408 =  n0323 & ~n0325;
assign n4409 =  n4407 & ~n4408;
assign n4410 =  n0324 & ~n0325;
assign n4411 =  n4409 & ~n4410;
assign n4412 =  n0081 & ~n0325;
assign n4413 =  n4411 & ~n4412;
assign n4414 =  n0078 & ~n0325;
assign n4415 =  n4413 & ~n4414;
assign n4416 =  n0072 & ~n0325;
assign n4417 =  n4415 & ~n4416;
assign n4418 =  n0066 & ~n0325;
assign n4419 =  n4417 & ~n4418;
assign n4420 =  n0042 & ~n0325;
assign n4421 =  n4419 & ~n4420;
assign n4422 =  n0041 & ~n0325;
assign n4423 =  n4421 & ~n4422;
assign n4424 =  n0036 & ~n0325;
assign n4425 =  n4423 & ~n4424;
assign n4426 = ~n0016 &  n0043;
assign n4427 = ~n0324 &  n4426;
assign n4428 =  n4425 & ~n4427;
assign n4429 =  n0016 &  n0048;
assign n4430 = ~n0323 &  n4429;
assign n4431 =  n4428 & ~n4430;
assign n4432 =  n0016 &  n0047;
assign n4433 = ~n0322 &  n4432;
assign n4434 =  n4431 & ~n4433;
assign n4435 = ~n0016 &  n0045;
assign n4436 = ~n0321 &  n4435;
assign n4437 =  n4434 & ~n4436;
assign n4438 =  n0015 &  n0020;
assign n4439 = ~n0320 &  n4438;
assign n4440 =  n4437 & ~n4439;
assign n4441 = ~n0015 &  n0018;
assign n4442 = ~n0319 &  n4441;
assign n4443 =  n4440 & ~n4442;
assign n4444 = ~n0015 &  n0044;
assign n4445 = ~n0318 &  n4444;
assign n4446 =  n4443 & ~n4445;
assign n4447 =  n0015 &  n0046;
assign n4448 = ~n0317 &  n4447;
assign n4449 =  n4446 & ~n4448;
assign n4450 =  n0308 & ~n0316;
assign n4451 =  n4449 & ~n4450;
assign n4452 =  n0309 & ~n0316;
assign n4453 =  n4451 & ~n4452;
assign n4454 =  n0310 & ~n0316;
assign n4455 =  n4453 & ~n4454;
assign n4456 =  n0311 & ~n0316;
assign n4457 =  n4455 & ~n4456;
assign n4458 =  n0312 & ~n0316;
assign n4459 =  n4457 & ~n4458;
assign n4460 =  n0313 & ~n0316;
assign n4461 =  n4459 & ~n4460;
assign n4462 =  n0314 & ~n0316;
assign n4463 =  n4461 & ~n4462;
assign n4464 =  n0080 & ~n0316;
assign n4465 =  n4463 & ~n4464;
assign n4466 =  n0077 & ~n0316;
assign n4467 =  n4465 & ~n4466;
assign n4468 =  n0071 & ~n0316;
assign n4469 =  n4467 & ~n4468;
assign n4470 =  n0063 & ~n0316;
assign n4471 =  n4469 & ~n4470;
assign n4472 =  n0315 & ~n0316;
assign n4473 =  n4471 & ~n4472;
assign n4474 =  n0029 & ~n0316;
assign n4475 =  n4473 & ~n4474;
assign n4476 =  n0028 & ~n0316;
assign n4477 =  n4475 & ~n4476;
assign n4478 =  n0023 & ~n0316;
assign n4479 =  n4477 & ~n4478;
assign n4480 =  n0015 &  n0033;
assign n4481 = ~n0315 &  n4480;
assign n4482 =  n4479 & ~n4481;
assign n4483 = ~n0016 &  n0030;
assign n4484 = ~n0314 &  n4483;
assign n4485 =  n4482 & ~n4484;
assign n4486 =  n0016 &  n0034;
assign n4487 = ~n0313 &  n4486;
assign n4488 =  n4485 & ~n4487;
assign n4489 =  n0016 &  n0035;
assign n4490 = ~n0312 &  n4489;
assign n4491 =  n4488 & ~n4490;
assign n4492 = ~n0016 &  n0032;
assign n4493 = ~n0311 &  n4492;
assign n4494 =  n4491 & ~n4493;
assign n4495 =  n0015 &  n0021;
assign n4496 = ~n0310 &  n4495;
assign n4497 =  n4494 & ~n4496;
assign n4498 = ~n0015 &  n0017;
assign n4499 = ~n0309 &  n4498;
assign n4500 =  n4497 & ~n4499;
assign n4501 = ~n0015 &  n0031;
assign n4502 = ~n0308 &  n4501;
assign n4503 =  n4500 & ~n4502;
assign n4504 =  n0302 &  n0898;
assign n4505 = ~n0307 &  n4504;
assign n4506 =  n4503 & ~n4505;
assign n4507 =  n0014 & ~n0306;
assign n4508 =  n4506 & ~n4507;
assign n4509 =  n0013 & ~n0306;
assign n4510 =  n4508 & ~n4509;
assign n4511 =  n0010 & ~n0305;
assign n4512 =  n4510 & ~n4511;
assign n4513 =  n0009 & ~n0305;
assign n4514 =  n4512 & ~n4513;
assign n4515 =  n0012 & ~n0304;
assign n4516 =  n4514 & ~n4515;
assign n4517 =  n0011 & ~n0304;
assign n4518 =  n4516 & ~n4517;
assign n4519 =  n0016 & ~n0303;
assign n4520 =  n4518 & ~n4519;
assign n4521 =  n0015 & ~n0303;
assign n4522 =  n4520 & ~n4521;
assign n4523 =  n0115 & ~n0302;
assign n4524 =  n4522 & ~n4523;
assign n4525 =  n0264 & ~n0302;
assign n4526 =  n4524 & ~n4525;
assign n4527 =  n0283 & ~n0302;
assign n4528 =  n4526 & ~n4527;
assign n4529 =  n0301 & ~n0302;
assign n4530 =  n4528 & ~n4529;
assign n4531 =  n0286 &  n0300;
assign n4532 = ~n0301 &  n4531;
assign n4533 =  n4530 & ~n4532;
assign n4534 =  n0287 & ~n0300;
assign n4535 =  n4533 & ~n4534;
assign n4536 =  n0288 & ~n0300;
assign n4537 =  n4535 & ~n4536;
assign n4538 =  n0293 & ~n0300;
assign n4539 =  n4537 & ~n4538;
assign n4540 =  n0298 & ~n0300;
assign n4541 =  n4539 & ~n4540;
assign n4542 =  n0299 & ~n0300;
assign n4543 =  n4541 & ~n4542;
assign n4544 =  n0249 &  n0912;
assign n4545 = ~n0299 &  n4544;
assign n4546 =  n4543 & ~n4545;
assign n4547 =  n0258 &  n2170;
assign n4548 = ~n0298 &  n4547;
assign n4549 =  n4546 & ~n4548;
assign n4550 =  n0294 & ~n0297;
assign n4551 =  n4549 & ~n4550;
assign n4552 =  n0295 & ~n0297;
assign n4553 =  n4551 & ~n4552;
assign n4554 =  n0296 & ~n0297;
assign n4555 =  n4553 & ~n4554;
assign n4556 = ~n0296 &  n2246;
assign n4557 =  n4555 & ~n4556;
assign n4558 =  n0215 &  n1780;
assign n4559 = ~n0295 &  n4558;
assign n4560 =  n4557 & ~n4559;
assign n4561 =  n0192 &  n4544;
assign n4562 = ~n0294 &  n4561;
assign n4563 =  n4560 & ~n4562;
assign n4564 =  n0292 &  n0912;
assign n4565 =  n0241 &  n4564;
assign n4566 = ~n0293 &  n4565;
assign n4567 =  n4563 & ~n4566;
assign n4568 =  n0289 & ~n0292;
assign n4569 =  n4567 & ~n4568;
assign n4570 =  n0290 & ~n0292;
assign n4571 =  n4569 & ~n4570;
assign n4572 =  n0291 & ~n0292;
assign n4573 =  n4571 & ~n4572;
assign n4574 = ~n0291 &  n2214;
assign n4575 =  n4573 & ~n4574;
assign n4576 =  n0232 &  n2246;
assign n4577 = ~n0290 &  n4576;
assign n4578 =  n4575 & ~n4577;
assign n4579 =  n0159 &  n4544;
assign n4580 = ~n0289 &  n4579;
assign n4581 =  n4578 & ~n4580;
assign n4582 =  n0258 &  n2246;
assign n4583 = ~n0288 &  n4582;
assign n4584 =  n4581 & ~n4583;
assign n4585 =  n0241 &  n2214;
assign n4586 = ~n0287 &  n4585;
assign n4587 =  n4584 & ~n4586;
assign n4588 =  n0160 & ~n0286;
assign n4589 =  n4587 & ~n4588;
assign n4590 =  n0193 & ~n0286;
assign n4591 =  n4589 & ~n4590;
assign n4592 =  n0284 & ~n0286;
assign n4593 =  n4591 & ~n4592;
assign n4594 =  n0285 & ~n0286;
assign n4595 =  n4593 & ~n4594;
assign n4596 =  n0198 & ~n0286;
assign n4597 =  n4595 & ~n4596;
assign n4598 =  n0228 &  n0912;
assign n4599 =  n0176 &  n4598;
assign n4600 = ~n0285 &  n4599;
assign n4601 =  n4597 & ~n4600;
assign n4602 =  n0266 &  n0912;
assign n4603 =  n0143 &  n4602;
assign n4604 = ~n0284 &  n4603;
assign n4605 =  n4601 & ~n4604;
assign n4606 =  n0268 &  n0282;
assign n4607 = ~n0283 &  n4606;
assign n4608 =  n4605 & ~n4607;
assign n4609 =  n0273 & ~n0282;
assign n4610 =  n4608 & ~n4609;
assign n4611 =  n0278 & ~n0282;
assign n4612 =  n4610 & ~n4611;
assign n4613 =  n0279 & ~n0282;
assign n4614 =  n4612 & ~n4613;
assign n4615 =  n0280 & ~n0282;
assign n4616 =  n4614 & ~n4615;
assign n4617 =  n0281 & ~n0282;
assign n4618 =  n4616 & ~n4617;
assign n4619 =  n0258 &  n0912;
assign n4620 = ~n0281 &  n4619;
assign n4621 =  n4618 & ~n4620;
assign n4622 =  n0176 &  n4544;
assign n4623 = ~n0280 &  n4622;
assign n4624 =  n4621 & ~n4623;
assign n4625 =  n0232 &  n0912;
assign n4626 =  n0241 &  n4625;
assign n4627 = ~n0279 &  n4626;
assign n4628 =  n4624 & ~n4627;
assign n4629 =  n0277 &  n4544;
assign n4630 = ~n0278 &  n4629;
assign n4631 =  n4628 & ~n4630;
assign n4632 =  n0274 & ~n0277;
assign n4633 =  n4631 & ~n4632;
assign n4634 =  n0275 & ~n0277;
assign n4635 =  n4633 & ~n4634;
assign n4636 =  n0276 & ~n0277;
assign n4637 =  n4635 & ~n4636;
assign n4638 = ~n0276 &  n2194;
assign n4639 =  n4637 & ~n4638;
assign n4640 =  n0143 &  n4625;
assign n4641 = ~n0275 &  n4640;
assign n4642 =  n4639 & ~n4641;
assign n4643 =  n0197 &  n4619;
assign n4644 = ~n0274 &  n4643;
assign n4645 =  n4642 & ~n4644;
assign n4646 =  n0241 &  n0912;
assign n4647 =  n0272 &  n4646;
assign n4648 = ~n0273 &  n4647;
assign n4649 =  n4645 & ~n4648;
assign n4650 =  n0269 & ~n0272;
assign n4651 =  n4649 & ~n4650;
assign n4652 =  n0270 & ~n0272;
assign n4653 =  n4651 & ~n4652;
assign n4654 =  n0271 & ~n0272;
assign n4655 =  n4653 & ~n4654;
assign n4656 = ~n0271 &  n4625;
assign n4657 =  n4655 & ~n4656;
assign n4658 =  n0176 &  n2214;
assign n4659 = ~n0270 &  n4658;
assign n4660 =  n4657 & ~n4659;
assign n4661 =  n0159 &  n4619;
assign n4662 = ~n0269 &  n4661;
assign n4663 =  n4660 & ~n4662;
assign n4664 =  n0265 & ~n0268;
assign n4665 =  n4663 & ~n4664;
assign n4666 =  n0267 & ~n0268;
assign n4667 =  n4665 & ~n4666;
assign n4668 =  n0221 & ~n0268;
assign n4669 =  n4667 & ~n4668;
assign n4670 =  n0226 & ~n0268;
assign n4671 =  n4669 & ~n4670;
assign n4672 =  n0227 & ~n0268;
assign n4673 =  n4671 & ~n4672;
assign n4674 =  n0266 &  n1780;
assign n4675 = ~n0267 &  n4674;
assign n4676 =  n4673 & ~n4675;
assign n4677 =  n0234 & ~n0266;
assign n4678 =  n4676 & ~n4677;
assign n4679 =  n0235 & ~n0266;
assign n4680 =  n4678 & ~n4679;
assign n4681 =  n0236 & ~n0266;
assign n4682 =  n4680 & ~n4681;
assign n4683 =  n0199 &  n2246;
assign n4684 = ~n0265 &  n4683;
assign n4685 =  n4682 & ~n4684;
assign n4686 =  n0237 &  n0263;
assign n4687 = ~n0264 &  n4686;
assign n4688 =  n4685 & ~n4687;
assign n4689 =  n0250 & ~n0263;
assign n4690 =  n4688 & ~n4689;
assign n4691 =  n0259 & ~n0263;
assign n4692 =  n4690 & ~n4691;
assign n4693 =  n0260 & ~n0263;
assign n4694 =  n4692 & ~n4693;
assign n4695 =  n0261 & ~n0263;
assign n4696 =  n4694 & ~n4695;
assign n4697 =  n0262 & ~n0263;
assign n4698 =  n4696 & ~n4697;
assign n4699 = ~n0262 &  n4646;
assign n4700 =  n4698 & ~n4699;
assign n4701 =  n0143 &  n4544;
assign n4702 = ~n0261 &  n4701;
assign n4703 =  n4700 & ~n4702;
assign n4704 =  n0258 &  n1780;
assign n4705 = ~n0260 &  n4704;
assign n4706 =  n4703 & ~n4705;
assign n4707 =  n0254 &  n4619;
assign n4708 = ~n0259 &  n4707;
assign n4709 =  n4706 & ~n4708;
assign n4710 =  n0255 & ~n0258;
assign n4711 =  n4709 & ~n4710;
assign n4712 =  n0256 & ~n0258;
assign n4713 =  n4711 & ~n4712;
assign n4714 =  n0257 & ~n0258;
assign n4715 =  n4713 & ~n4714;
assign n4716 = ~n0069 &  n0923;
assign n4717 = ~n0068 &  n4716;
assign n4718 = ~n0073 &  n4717;
assign n4719 = ~n0082 &  n4718;
assign n4720 =  n0174 &  n4719;
assign n4721 =  n0173 &  n4720;
assign n4722 =  n0107 &  n4721;
assign n4723 =  n0172 &  n4722;
assign n4724 =  n0106 &  n4723;
assign n4725 =  n0105 &  n4724;
assign n4726 =  n0103 &  n4725;
assign n4727 =  n0171 &  n4726;
assign n4728 = ~n0257 &  n4727;
assign n4729 =  n4715 & ~n4728;
assign n4730 = ~n0066 & ~n0081;
assign n4731 = ~n0040 &  n4730;
assign n4732 = ~n0065 &  n4731;
assign n4733 = ~n0072 &  n4732;
assign n4734 = ~n0042 &  n4733;
assign n4735 =  n0099 &  n4734;
assign n4736 = ~n0041 &  n4735;
assign n4737 =  n0097 &  n4736;
assign n4738 =  n0169 &  n4737;
assign n4739 =  n0168 &  n4738;
assign n4740 =  n0167 &  n4739;
assign n4741 =  n0095 &  n4740;
assign n4742 =  n0094 &  n4741;
assign n4743 =  n0166 &  n4742;
assign n4744 = ~n0256 &  n4743;
assign n4745 =  n4729 & ~n4744;
assign n4746 = ~n0028 & ~n0029;
assign n4747 = ~n0027 &  n4746;
assign n4748 = ~n0063 &  n4747;
assign n4749 = ~n0062 &  n4748;
assign n4750 = ~n0071 &  n4749;
assign n4751 = ~n0080 &  n4750;
assign n4752 =  n0089 &  n4751;
assign n4753 =  n0164 &  n4752;
assign n4754 =  n0163 &  n4753;
assign n4755 =  n0088 &  n4754;
assign n4756 =  n0085 &  n4755;
assign n4757 =  n0084 &  n4756;
assign n4758 =  n0162 &  n4757;
assign n4759 =  n0161 &  n4758;
assign n4760 = ~n0255 &  n4759;
assign n4761 =  n4745 & ~n4760;
assign n4762 =  n0251 & ~n0254;
assign n4763 =  n4761 & ~n4762;
assign n4764 =  n0252 & ~n0254;
assign n4765 =  n4763 & ~n4764;
assign n4766 =  n0253 & ~n0254;
assign n4767 =  n4765 & ~n4766;
assign n4768 = ~n0253 &  n1780;
assign n4769 =  n4767 & ~n4768;
assign n4770 =  n0143 &  n2246;
assign n4771 = ~n0252 &  n4770;
assign n4772 =  n4769 & ~n4771;
assign n4773 =  n0241 &  n1784;
assign n4774 = ~n0251 &  n4773;
assign n4775 =  n4772 & ~n4774;
assign n4776 =  n0245 &  n4544;
assign n4777 = ~n0250 &  n4776;
assign n4778 =  n4775 & ~n4777;
assign n4779 =  n0246 & ~n0249;
assign n4780 =  n4778 & ~n4779;
assign n4781 =  n0247 & ~n0249;
assign n4782 =  n4780 & ~n4781;
assign n4783 =  n0248 & ~n0249;
assign n4784 =  n4782 & ~n4783;
assign n4785 = ~n0068 &  n0923;
assign n4786 = ~n0051 &  n4785;
assign n4787 = ~n0073 &  n4786;
assign n4788 = ~n0082 &  n4787;
assign n4789 =  n0213 &  n4788;
assign n4790 =  n0212 &  n4789;
assign n4791 =  n0107 &  n4790;
assign n4792 =  n0211 &  n4791;
assign n4793 =  n0106 &  n4792;
assign n4794 =  n0105 &  n4793;
assign n4795 =  n0103 &  n4794;
assign n4796 =  n0210 &  n4795;
assign n4797 = ~n0248 &  n4796;
assign n4798 =  n4784 & ~n4797;
assign n4799 = ~n0038 & ~n0081;
assign n4800 = ~n0040 &  n4799;
assign n4801 = ~n0065 &  n4800;
assign n4802 = ~n0072 &  n4801;
assign n4803 = ~n0042 &  n4802;
assign n4804 =  n0099 &  n4803;
assign n4805 = ~n0041 &  n4804;
assign n4806 =  n0097 &  n4805;
assign n4807 =  n0208 &  n4806;
assign n4808 =  n0095 &  n4807;
assign n4809 =  n0094 &  n4808;
assign n4810 =  n0207 &  n4809;
assign n4811 =  n0206 &  n4810;
assign n4812 =  n0205 &  n4811;
assign n4813 = ~n0247 &  n4812;
assign n4814 =  n4798 & ~n4813;
assign n4815 = ~n0025 & ~n0028;
assign n4816 = ~n0029 &  n4815;
assign n4817 = ~n0027 &  n4816;
assign n4818 =  n0203 &  n4817;
assign n4819 = ~n0062 &  n4818;
assign n4820 = ~n0071 &  n4819;
assign n4821 = ~n0080 &  n4820;
assign n4822 =  n0089 &  n4821;
assign n4823 =  n0088 &  n4822;
assign n4824 =  n0085 &  n4823;
assign n4825 =  n0084 &  n4824;
assign n4826 =  n0202 &  n4825;
assign n4827 =  n0201 &  n4826;
assign n4828 =  n0200 &  n4827;
assign n4829 = ~n0246 &  n4828;
assign n4830 =  n4814 & ~n4829;
assign n4831 =  n0242 & ~n0245;
assign n4832 =  n4830 & ~n4831;
assign n4833 =  n0243 & ~n0245;
assign n4834 =  n4832 & ~n4833;
assign n4835 =  n0244 & ~n0245;
assign n4836 =  n4834 & ~n4835;
assign n4837 = ~n0244 &  n1878;
assign n4838 =  n4836 & ~n4837;
assign n4839 =  n0176 &  n1780;
assign n4840 = ~n0243 &  n4839;
assign n4841 =  n4838 & ~n4840;
assign n4842 =  n0197 &  n4646;
assign n4843 = ~n0242 &  n4842;
assign n4844 =  n4841 & ~n4843;
assign n4845 =  n0238 & ~n0241;
assign n4846 =  n4844 & ~n4845;
assign n4847 =  n0239 & ~n0241;
assign n4848 =  n4846 & ~n4847;
assign n4849 =  n0240 & ~n0241;
assign n4850 =  n4848 & ~n4849;
assign n4851 = ~n0076 &  n0922;
assign n4852 = ~n0069 &  n4851;
assign n4853 = ~n0068 &  n4852;
assign n4854 = ~n0073 &  n4853;
assign n4855 = ~n0082 &  n4854;
assign n4856 =  n0107 &  n4855;
assign n4857 =  n0141 &  n4856;
assign n4858 =  n0106 &  n4857;
assign n4859 =  n0105 &  n4858;
assign n4860 =  n0103 &  n4859;
assign n4861 =  n0139 &  n4860;
assign n4862 =  n0136 &  n4861;
assign n4863 =  n0135 &  n4862;
assign n4864 = ~n0240 &  n4863;
assign n4865 =  n4850 & ~n4864;
assign n4866 = ~n0075 &  n4732;
assign n4867 = ~n0072 &  n4866;
assign n4868 =  n0099 &  n4867;
assign n4869 = ~n0041 &  n4868;
assign n4870 =  n0097 &  n4869;
assign n4871 =  n0095 &  n4870;
assign n4872 =  n0094 &  n4871;
assign n4873 =  n0130 &  n4872;
assign n4874 =  n0128 &  n4873;
assign n4875 =  n0126 &  n4874;
assign n4876 =  n0125 &  n4875;
assign n4877 = ~n0239 &  n4876;
assign n4878 =  n4865 & ~n4877;
assign n4879 = ~n0027 & ~n0028;
assign n4880 = ~n0063 &  n4879;
assign n4881 = ~n0062 &  n4880;
assign n4882 = ~n0074 &  n4881;
assign n4883 = ~n0071 &  n4882;
assign n4884 = ~n0080 &  n4883;
assign n4885 =  n0089 &  n4884;
assign n4886 =  n0122 &  n4885;
assign n4887 =  n0088 &  n4886;
assign n4888 =  n0085 &  n4887;
assign n4889 =  n0084 &  n4888;
assign n4890 =  n0119 &  n4889;
assign n4891 =  n0118 &  n4890;
assign n4892 =  n0117 &  n4891;
assign n4893 = ~n0238 &  n4892;
assign n4894 =  n4878 & ~n4893;
assign n4895 =  n0216 & ~n0237;
assign n4896 =  n4894 & ~n4895;
assign n4897 =  n0233 & ~n0237;
assign n4898 =  n4896 & ~n4897;
assign n4899 =  n0234 & ~n0237;
assign n4900 =  n4898 & ~n4899;
assign n4901 =  n0235 & ~n0237;
assign n4902 =  n4900 & ~n4901;
assign n4903 =  n0236 & ~n0237;
assign n4904 =  n4902 & ~n4903;
assign n4905 = ~n0236 &  n2174;
assign n4906 =  n4904 & ~n4905;
assign n4907 =  n0197 &  n2214;
assign n4908 = ~n0235 &  n4907;
assign n4909 =  n4906 & ~n4908;
assign n4910 =  n0232 &  n1784;
assign n4911 = ~n0234 &  n4910;
assign n4912 =  n4909 & ~n4911;
assign n4913 =  n0228 &  n4625;
assign n4914 = ~n0233 &  n4913;
assign n4915 =  n4912 & ~n4914;
assign n4916 =  n0229 & ~n0232;
assign n4917 =  n4915 & ~n4916;
assign n4918 =  n0230 & ~n0232;
assign n4919 =  n4917 & ~n4918;
assign n4920 =  n0231 & ~n0232;
assign n4921 =  n4919 & ~n4920;
assign n4922 = ~n0076 &  n2260;
assign n4923 = ~n0052 &  n4922;
assign n4924 = ~n0069 &  n4923;
assign n4925 = ~n0068 &  n4924;
assign n4926 = ~n0073 &  n4925;
assign n4927 =  n0174 &  n4926;
assign n4928 =  n0173 &  n4927;
assign n4929 =  n0156 &  n4928;
assign n4930 =  n0155 &  n4929;
assign n4931 =  n0172 &  n4930;
assign n4932 =  n0154 &  n4931;
assign n4933 =  n0171 &  n4932;
assign n4934 = ~n0231 &  n4933;
assign n4935 =  n4921 & ~n4934;
assign n4936 = ~n0066 &  n2275;
assign n4937 = ~n0040 &  n4936;
assign n4938 = ~n0065 &  n4937;
assign n4939 = ~n0075 &  n4938;
assign n4940 = ~n0072 &  n4939;
assign n4941 = ~n0041 &  n4940;
assign n4942 =  n0151 &  n4941;
assign n4943 =  n0169 &  n4942;
assign n4944 =  n0168 &  n4943;
assign n4945 =  n0150 &  n4944;
assign n4946 =  n0167 &  n4945;
assign n4947 =  n0149 &  n4946;
assign n4948 =  n0166 &  n4947;
assign n4949 = ~n0230 &  n4948;
assign n4950 =  n4935 & ~n4949;
assign n4951 = ~n0026 &  n4879;
assign n4952 = ~n0063 &  n4951;
assign n4953 = ~n0062 &  n4952;
assign n4954 = ~n0074 &  n4953;
assign n4955 = ~n0071 &  n4954;
assign n4956 =  n0147 &  n4955;
assign n4957 =  n0146 &  n4956;
assign n4958 =  n0145 &  n4957;
assign n4959 =  n0164 &  n4958;
assign n4960 =  n0163 &  n4959;
assign n4961 =  n0144 &  n4960;
assign n4962 =  n0162 &  n4961;
assign n4963 =  n0161 &  n4962;
assign n4964 = ~n0229 &  n4963;
assign n4965 =  n4950 & ~n4964;
assign n4966 =  n0221 & ~n0228;
assign n4967 =  n4965 & ~n4966;
assign n4968 =  n0226 & ~n0228;
assign n4969 =  n4967 & ~n4968;
assign n4970 =  n0227 & ~n0228;
assign n4971 =  n4969 & ~n4970;
assign n4972 = ~n0227 &  n1784;
assign n4973 =  n4971 & ~n4972;
assign n4974 =  n0197 &  n2246;
assign n4975 = ~n0226 &  n4974;
assign n4976 =  n4973 & ~n4975;
assign n4977 =  n0222 & ~n0225;
assign n4978 =  n4976 & ~n4977;
assign n4979 =  n0223 & ~n0225;
assign n4980 =  n4978 & ~n4979;
assign n4981 =  n0224 & ~n0225;
assign n4982 =  n4980 & ~n4981;
assign n4983 = ~n0052 &  n4851;
assign n4984 = ~n0068 &  n4983;
assign n4985 = ~n0051 &  n4984;
assign n4986 = ~n0073 &  n4985;
assign n4987 =  n0190 &  n4986;
assign n4988 =  n0213 &  n4987;
assign n4989 =  n0212 &  n4988;
assign n4990 =  n0189 &  n4989;
assign n4991 =  n0188 &  n4990;
assign n4992 =  n0211 &  n4991;
assign n4993 =  n0210 &  n4992;
assign n4994 =  n0187 &  n4993;
assign n4995 = ~n0224 &  n4994;
assign n4996 =  n4982 & ~n4995;
assign n4997 = ~n0040 &  n0938;
assign n4998 = ~n0065 &  n4997;
assign n4999 = ~n0075 &  n4998;
assign n5000 = ~n0072 &  n4999;
assign n5001 = ~n0041 &  n5000;
assign n5002 =  n0185 &  n5001;
assign n5003 =  n0184 &  n5002;
assign n5004 =  n0183 &  n5003;
assign n5005 =  n0208 &  n5004;
assign n5006 =  n0182 &  n5005;
assign n5007 =  n0207 &  n5006;
assign n5008 =  n0206 &  n5007;
assign n5009 =  n0205 &  n5008;
assign n5010 = ~n0223 &  n5009;
assign n5011 =  n4996 & ~n5010;
assign n5012 = ~n0027 &  n4815;
assign n5013 = ~n0026 &  n5012;
assign n5014 =  n0203 &  n5013;
assign n5015 = ~n0062 &  n5014;
assign n5016 = ~n0074 &  n5015;
assign n5017 = ~n0071 &  n5016;
assign n5018 =  n0180 &  n5017;
assign n5019 =  n0179 &  n5018;
assign n5020 =  n0178 &  n5019;
assign n5021 =  n0202 &  n5020;
assign n5022 =  n0201 &  n5021;
assign n5023 =  n0200 &  n5022;
assign n5024 =  n0177 &  n5023;
assign n5025 = ~n0222 &  n5024;
assign n5026 =  n5011 & ~n5025;
assign n5027 =  n0159 &  n1780;
assign n5028 = ~n0221 &  n5027;
assign n5029 =  n5026 & ~n5028;
assign n5030 =  n0217 & ~n0220;
assign n5031 =  n5029 & ~n5030;
assign n5032 =  n0218 & ~n0220;
assign n5033 =  n5031 & ~n5032;
assign n5034 =  n0219 & ~n0220;
assign n5035 =  n5033 & ~n5034;
assign n5036 = ~n0053 & ~n0055;
assign n5037 = ~n0052 &  n5036;
assign n5038 = ~n0069 &  n5037;
assign n5039 = ~n0068 &  n5038;
assign n5040 = ~n0073 &  n5039;
assign n5041 = ~n0070 &  n5040;
assign n5042 =  n0190 &  n5041;
assign n5043 =  n0189 &  n5042;
assign n5044 =  n0141 &  n5043;
assign n5045 =  n0188 &  n5044;
assign n5046 =  n0139 &  n5045;
assign n5047 =  n0136 &  n5046;
assign n5048 =  n0187 &  n5047;
assign n5049 =  n0135 &  n5048;
assign n5050 = ~n0219 &  n5049;
assign n5051 =  n5035 & ~n5050;
assign n5052 = ~n0039 & ~n0067;
assign n5053 = ~n0066 &  n5052;
assign n5054 = ~n0040 &  n5053;
assign n5055 = ~n0065 &  n5054;
assign n5056 = ~n0072 &  n5055;
assign n5057 = ~n0042 &  n5056;
assign n5058 =  n0185 &  n5057;
assign n5059 =  n0184 &  n5058;
assign n5060 =  n0183 &  n5059;
assign n5061 =  n0182 &  n5060;
assign n5062 =  n0130 &  n5061;
assign n5063 =  n0128 &  n5062;
assign n5064 =  n0126 &  n5063;
assign n5065 =  n0125 &  n5064;
assign n5066 = ~n0218 &  n5065;
assign n5067 =  n5051 & ~n5066;
assign n5068 = ~n0027 & ~n0029;
assign n5069 = ~n0026 &  n5068;
assign n5070 = ~n0064 &  n5069;
assign n5071 = ~n0063 &  n5070;
assign n5072 = ~n0062 &  n5071;
assign n5073 = ~n0071 &  n5072;
assign n5074 =  n0180 &  n5073;
assign n5075 =  n0122 &  n5074;
assign n5076 =  n0179 &  n5075;
assign n5077 =  n0178 &  n5076;
assign n5078 =  n0177 &  n5077;
assign n5079 =  n0119 &  n5078;
assign n5080 =  n0118 &  n5079;
assign n5081 =  n0117 &  n5080;
assign n5082 = ~n0217 &  n5081;
assign n5083 =  n5067 & ~n5082;
assign n5084 =  n0199 &  n2214;
assign n5085 = ~n0216 &  n5084;
assign n5086 =  n5083 & ~n5085;
assign n5087 =  n0204 & ~n0215;
assign n5088 =  n5086 & ~n5087;
assign n5089 =  n0209 & ~n0215;
assign n5090 =  n5088 & ~n5089;
assign n5091 =  n0214 & ~n0215;
assign n5092 =  n5090 & ~n5091;
assign n5093 = ~n0068 &  n2262;
assign n5094 = ~n0051 &  n5093;
assign n5095 = ~n0073 &  n5094;
assign n5096 =  n0213 &  n5095;
assign n5097 =  n0156 &  n5096;
assign n5098 =  n0212 &  n5097;
assign n5099 =  n0155 &  n5098;
assign n5100 =  n0211 &  n5099;
assign n5101 =  n0210 &  n5100;
assign n5102 =  n0154 &  n5101;
assign n5103 = ~n0214 &  n5102;
assign n5104 =  n5092 & ~n5103;
assign n5105 = ~n0061 & ~n0213;
assign n5106 =  n5104 & ~n5105;
assign n5107 = ~n0010 & ~n0213;
assign n5108 =  n5106 & ~n5107;
assign n5109 = ~n0057 & ~n0212;
assign n5110 =  n5108 & ~n5109;
assign n5111 =  n0009 & ~n0212;
assign n5112 =  n5110 & ~n5111;
assign n5113 = ~n0059 & ~n0211;
assign n5114 =  n5112 & ~n5113;
assign n5115 = ~n0009 & ~n0211;
assign n5116 =  n5114 & ~n5115;
assign n5117 = ~n0058 & ~n0210;
assign n5118 =  n5116 & ~n5117;
assign n5119 =  n0010 & ~n0210;
assign n5120 =  n5118 & ~n5119;
assign n5121 = ~n0038 &  n2275;
assign n5122 = ~n0040 &  n5121;
assign n5123 = ~n0065 &  n5122;
assign n5124 = ~n0072 &  n5123;
assign n5125 = ~n0042 &  n5124;
assign n5126 = ~n0041 &  n5125;
assign n5127 =  n0151 &  n5126;
assign n5128 =  n0208 &  n5127;
assign n5129 =  n0150 &  n5128;
assign n5130 =  n0149 &  n5129;
assign n5131 =  n0207 &  n5130;
assign n5132 =  n0206 &  n5131;
assign n5133 =  n0205 &  n5132;
assign n5134 = ~n0209 &  n5133;
assign n5135 =  n5120 & ~n5134;
assign n5136 = ~n0044 & ~n0208;
assign n5137 =  n5135 & ~n5136;
assign n5138 =  n0009 & ~n0208;
assign n5139 =  n5137 & ~n5138;
assign n5140 = ~n0046 & ~n0207;
assign n5141 =  n5139 & ~n5140;
assign n5142 = ~n0009 & ~n0207;
assign n5143 =  n5141 & ~n5142;
assign n5144 = ~n0048 & ~n0206;
assign n5145 =  n5143 & ~n5144;
assign n5146 = ~n0010 & ~n0206;
assign n5147 =  n5145 & ~n5146;
assign n5148 = ~n0045 & ~n0205;
assign n5149 =  n5147 & ~n5148;
assign n5150 =  n0010 & ~n0205;
assign n5151 =  n5149 & ~n5150;
assign n5152 = ~n0026 &  n4817;
assign n5153 =  n0203 &  n5152;
assign n5154 = ~n0062 &  n5153;
assign n5155 = ~n0071 &  n5154;
assign n5156 =  n0147 &  n5155;
assign n5157 =  n0146 &  n5156;
assign n5158 =  n0145 &  n5157;
assign n5159 =  n0202 &  n5158;
assign n5160 =  n0144 &  n5159;
assign n5161 =  n0201 &  n5160;
assign n5162 =  n0200 &  n5161;
assign n5163 = ~n0204 &  n5162;
assign n5164 =  n5151 & ~n5163;
assign n5165 = ~n0033 & ~n0203;
assign n5166 =  n5164 & ~n5165;
assign n5167 = ~n0009 & ~n0203;
assign n5168 =  n5166 & ~n5167;
assign n5169 = ~n0031 & ~n0202;
assign n5170 =  n5168 & ~n5169;
assign n5171 =  n0009 & ~n0202;
assign n5172 =  n5170 & ~n5171;
assign n5173 = ~n0035 & ~n0201;
assign n5174 =  n5172 & ~n5173;
assign n5175 = ~n0010 & ~n0201;
assign n5176 =  n5174 & ~n5175;
assign n5177 = ~n0032 & ~n0200;
assign n5178 =  n5176 & ~n5177;
assign n5179 =  n0010 & ~n0200;
assign n5180 =  n5178 & ~n5179;
assign n5181 =  n0160 & ~n0199;
assign n5182 =  n5180 & ~n5181;
assign n5183 =  n0193 & ~n0199;
assign n5184 =  n5182 & ~n5183;
assign n5185 =  n0198 & ~n0199;
assign n5186 =  n5184 & ~n5185;
assign n5187 = ~n0198 &  n1882;
assign n5188 =  n5186 & ~n5187;
assign n5189 =  n0194 & ~n0197;
assign n5190 =  n5188 & ~n5189;
assign n5191 =  n0195 & ~n0197;
assign n5192 =  n5190 & ~n5191;
assign n5193 =  n0196 & ~n0197;
assign n5194 =  n5192 & ~n5193;
assign n5195 = ~n0054 & ~n0055;
assign n5196 = ~n0052 &  n5195;
assign n5197 = ~n0050 &  n5196;
assign n5198 = ~n0069 &  n5197;
assign n5199 = ~n0068 &  n5198;
assign n5200 = ~n0079 &  n5199;
assign n5201 =  n0108 &  n5200;
assign n5202 =  n0140 &  n5201;
assign n5203 =  n0104 &  n5202;
assign n5204 =  n0102 &  n5203;
assign n5205 =  n0138 &  n5204;
assign n5206 =  n0137 &  n5205;
assign n5207 =  n0101 &  n5206;
assign n5208 =  n0134 &  n5207;
assign n5209 = ~n0196 &  n5208;
assign n5210 =  n5194 & ~n5209;
assign n5211 = ~n0037 & ~n0039;
assign n5212 = ~n0066 &  n5211;
assign n5213 = ~n0065 &  n5212;
assign n5214 = ~n0078 &  n5213;
assign n5215 = ~n0042 &  n5214;
assign n5216 = ~n0041 &  n5215;
assign n5217 =  n0098 &  n5216;
assign n5218 =  n0132 &  n5217;
assign n5219 =  n0096 &  n5218;
assign n5220 =  n0131 &  n5219;
assign n5221 =  n0093 &  n5220;
assign n5222 =  n0129 &  n5221;
assign n5223 =  n0127 &  n5222;
assign n5224 =  n0092 &  n5223;
assign n5225 = ~n0195 &  n5224;
assign n5226 =  n5210 & ~n5225;
assign n5227 = ~n0024 & ~n0028;
assign n5228 = ~n0029 &  n5227;
assign n5229 = ~n0026 &  n5228;
assign n5230 =  n0090 &  n5229;
assign n5231 = ~n0063 &  n5230;
assign n5232 = ~n0062 &  n5231;
assign n5233 = ~n0077 &  n5232;
assign n5234 =  n0123 &  n5233;
assign n5235 =  n0087 &  n5234;
assign n5236 =  n0086 &  n5235;
assign n5237 =  n0121 &  n5236;
assign n5238 =  n0083 &  n5237;
assign n5239 =  n0120 &  n5238;
assign n5240 =  n0116 &  n5239;
assign n5241 = ~n0194 &  n5240;
assign n5242 =  n5226 & ~n5241;
assign n5243 =  n0176 &  n1784;
assign n5244 = ~n0193 &  n5243;
assign n5245 =  n5242 & ~n5244;
assign n5246 =  n0181 & ~n0192;
assign n5247 =  n5245 & ~n5246;
assign n5248 =  n0186 & ~n0192;
assign n5249 =  n5247 & ~n5248;
assign n5250 =  n0191 & ~n0192;
assign n5251 =  n5249 & ~n5250;
assign n5252 = ~n0069 &  n5196;
assign n5253 = ~n0068 &  n5252;
assign n5254 = ~n0079 &  n5253;
assign n5255 = ~n0073 &  n5254;
assign n5256 =  n0190 &  n5255;
assign n5257 =  n0108 &  n5256;
assign n5258 =  n0189 &  n5257;
assign n5259 =  n0188 &  n5258;
assign n5260 =  n0104 &  n5259;
assign n5261 =  n0102 &  n5260;
assign n5262 =  n0187 &  n5261;
assign n5263 =  n0101 &  n5262;
assign n5264 = ~n0191 &  n5263;
assign n5265 =  n5251 & ~n5264;
assign n5266 = ~n0011 & ~n0190;
assign n5267 =  n5265 & ~n5266;
assign n5268 = ~n0022 & ~n0190;
assign n5269 =  n5267 & ~n5268;
assign n5270 = ~n0060 & ~n0189;
assign n5271 =  n5269 & ~n5270;
assign n5272 = ~n0012 & ~n0189;
assign n5273 =  n5271 & ~n5272;
assign n5274 = ~n0019 & ~n0188;
assign n5275 =  n5273 & ~n5274;
assign n5276 =  n0011 & ~n0188;
assign n5277 =  n5275 & ~n5276;
assign n5278 = ~n0056 & ~n0187;
assign n5279 =  n5277 & ~n5278;
assign n5280 =  n0012 & ~n0187;
assign n5281 =  n5279 & ~n5280;
assign n5282 = ~n0039 & ~n0066;
assign n5283 = ~n0065 &  n5282;
assign n5284 = ~n0078 &  n5283;
assign n5285 = ~n0072 &  n5284;
assign n5286 = ~n0042 &  n5285;
assign n5287 = ~n0041 &  n5286;
assign n5288 =  n0098 &  n5287;
assign n5289 =  n0185 &  n5288;
assign n5290 =  n0184 &  n5289;
assign n5291 =  n0183 &  n5290;
assign n5292 =  n0096 &  n5291;
assign n5293 =  n0182 &  n5292;
assign n5294 =  n0093 &  n5293;
assign n5295 =  n0092 &  n5294;
assign n5296 = ~n0186 &  n5295;
assign n5297 =  n5281 & ~n5296;
assign n5298 = ~n0011 & ~n0185;
assign n5299 =  n5297 & ~n5298;
assign n5300 = ~n0020 & ~n0185;
assign n5301 =  n5299 & ~n5300;
assign n5302 = ~n0047 & ~n0184;
assign n5303 =  n5301 & ~n5302;
assign n5304 = ~n0012 & ~n0184;
assign n5305 =  n5303 & ~n5304;
assign n5306 = ~n0043 & ~n0183;
assign n5307 =  n5305 & ~n5306;
assign n5308 =  n0012 & ~n0183;
assign n5309 =  n5307 & ~n5308;
assign n5310 = ~n0018 & ~n0182;
assign n5311 =  n5309 & ~n5310;
assign n5312 =  n0011 & ~n0182;
assign n5313 =  n5311 & ~n5312;
assign n5314 = ~n0026 &  n4746;
assign n5315 =  n0090 &  n5314;
assign n5316 = ~n0063 &  n5315;
assign n5317 = ~n0062 &  n5316;
assign n5318 = ~n0077 &  n5317;
assign n5319 = ~n0071 &  n5318;
assign n5320 =  n0180 &  n5319;
assign n5321 =  n0179 &  n5320;
assign n5322 =  n0087 &  n5321;
assign n5323 =  n0086 &  n5322;
assign n5324 =  n0178 &  n5323;
assign n5325 =  n0083 &  n5324;
assign n5326 =  n0177 &  n5325;
assign n5327 = ~n0181 &  n5326;
assign n5328 =  n5313 & ~n5327;
assign n5329 = ~n0011 & ~n0180;
assign n5330 =  n5328 & ~n5329;
assign n5331 = ~n0021 & ~n0180;
assign n5332 =  n5330 & ~n5331;
assign n5333 = ~n0017 & ~n0179;
assign n5334 =  n5332 & ~n5333;
assign n5335 =  n0011 & ~n0179;
assign n5336 =  n5334 & ~n5335;
assign n5337 = ~n0034 & ~n0178;
assign n5338 =  n5336 & ~n5337;
assign n5339 = ~n0012 & ~n0178;
assign n5340 =  n5338 & ~n5339;
assign n5341 = ~n0030 & ~n0177;
assign n5342 =  n5340 & ~n5341;
assign n5343 =  n0012 & ~n0177;
assign n5344 =  n5342 & ~n5343;
assign n5345 =  n0165 & ~n0176;
assign n5346 =  n5344 & ~n5345;
assign n5347 =  n0170 & ~n0176;
assign n5348 =  n5346 & ~n5347;
assign n5349 =  n0175 & ~n0176;
assign n5350 =  n5348 & ~n5349;
assign n5351 = ~n0050 &  n5037;
assign n5352 = ~n0069 &  n5351;
assign n5353 = ~n0068 &  n5352;
assign n5354 = ~n0070 &  n5353;
assign n5355 =  n0174 &  n5354;
assign n5356 =  n0173 &  n5355;
assign n5357 =  n0140 &  n5356;
assign n5358 =  n0172 &  n5357;
assign n5359 =  n0138 &  n5358;
assign n5360 =  n0137 &  n5359;
assign n5361 =  n0171 &  n5360;
assign n5362 =  n0134 &  n5361;
assign n5363 = ~n0175 &  n5362;
assign n5364 =  n5350 & ~n5363;
assign n5365 = ~n0061 & ~n0174;
assign n5366 =  n5364 & ~n5365;
assign n5367 = ~n0012 & ~n0174;
assign n5368 =  n5366 & ~n5367;
assign n5369 = ~n0059 & ~n0173;
assign n5370 =  n5368 & ~n5369;
assign n5371 = ~n0011 & ~n0173;
assign n5372 =  n5370 & ~n5371;
assign n5373 = ~n0057 & ~n0172;
assign n5374 =  n5372 & ~n5373;
assign n5375 =  n0011 & ~n0172;
assign n5376 =  n5374 & ~n5375;
assign n5377 = ~n0058 & ~n0171;
assign n5378 =  n5376 & ~n5377;
assign n5379 =  n0012 & ~n0171;
assign n5380 =  n5378 & ~n5379;
assign n5381 = ~n0067 &  n5211;
assign n5382 = ~n0066 &  n5381;
assign n5383 = ~n0040 &  n5382;
assign n5384 = ~n0065 &  n5383;
assign n5385 = ~n0042 &  n5384;
assign n5386 =  n0169 &  n5385;
assign n5387 =  n0168 &  n5386;
assign n5388 =  n0132 &  n5387;
assign n5389 =  n0167 &  n5388;
assign n5390 =  n0131 &  n5389;
assign n5391 =  n0129 &  n5390;
assign n5392 =  n0127 &  n5391;
assign n5393 =  n0166 &  n5392;
assign n5394 = ~n0170 &  n5393;
assign n5395 =  n5380 & ~n5394;
assign n5396 = ~n0048 & ~n0169;
assign n5397 =  n5395 & ~n5396;
assign n5398 = ~n0012 & ~n0169;
assign n5399 =  n5397 & ~n5398;
assign n5400 = ~n0044 & ~n0168;
assign n5401 =  n5399 & ~n5400;
assign n5402 =  n0011 & ~n0168;
assign n5403 =  n5401 & ~n5402;
assign n5404 = ~n0046 & ~n0167;
assign n5405 =  n5403 & ~n5404;
assign n5406 = ~n0011 & ~n0167;
assign n5407 =  n5405 & ~n5406;
assign n5408 = ~n0045 & ~n0166;
assign n5409 =  n5407 & ~n5408;
assign n5410 =  n0012 & ~n0166;
assign n5411 =  n5409 & ~n5410;
assign n5412 = ~n0024 & ~n0029;
assign n5413 = ~n0027 &  n5412;
assign n5414 = ~n0026 &  n5413;
assign n5415 = ~n0064 &  n5414;
assign n5416 = ~n0063 &  n5415;
assign n5417 = ~n0062 &  n5416;
assign n5418 =  n0123 &  n5417;
assign n5419 =  n0164 &  n5418;
assign n5420 =  n0163 &  n5419;
assign n5421 =  n0121 &  n5420;
assign n5422 =  n0120 &  n5421;
assign n5423 =  n0162 &  n5422;
assign n5424 =  n0161 &  n5423;
assign n5425 =  n0116 &  n5424;
assign n5426 = ~n0165 &  n5425;
assign n5427 =  n5411 & ~n5426;
assign n5428 = ~n0031 & ~n0164;
assign n5429 =  n5427 & ~n5428;
assign n5430 =  n0011 & ~n0164;
assign n5431 =  n5429 & ~n5430;
assign n5432 = ~n0033 & ~n0163;
assign n5433 =  n5431 & ~n5432;
assign n5434 = ~n0011 & ~n0163;
assign n5435 =  n5433 & ~n5434;
assign n5436 = ~n0035 & ~n0162;
assign n5437 =  n5435 & ~n5436;
assign n5438 = ~n0012 & ~n0162;
assign n5439 =  n5437 & ~n5438;
assign n5440 = ~n0032 & ~n0161;
assign n5441 =  n5439 & ~n5440;
assign n5442 =  n0012 & ~n0161;
assign n5443 =  n5441 & ~n5442;
assign n5444 =  n0143 &  n2174;
assign n5445 = ~n0160 &  n5444;
assign n5446 =  n5443 & ~n5445;
assign n5447 =  n0148 & ~n0159;
assign n5448 =  n5446 & ~n5447;
assign n5449 =  n0153 & ~n0159;
assign n5450 =  n5448 & ~n5449;
assign n5451 =  n0158 & ~n0159;
assign n5452 =  n5450 & ~n5451;
assign n5453 = ~n0055 &  n0157;
assign n5454 = ~n0052 &  n5453;
assign n5455 = ~n0069 &  n5454;
assign n5456 = ~n0068 &  n5455;
assign n5457 = ~n0079 &  n5456;
assign n5458 = ~n0073 &  n5457;
assign n5459 = ~n0070 &  n5458;
assign n5460 =  n0108 &  n5459;
assign n5461 =  n0156 &  n5460;
assign n5462 =  n0155 &  n5461;
assign n5463 =  n0104 &  n5462;
assign n5464 =  n0102 &  n5463;
assign n5465 =  n0154 &  n5464;
assign n5466 =  n0101 &  n5465;
assign n5467 = ~n0158 &  n5466;
assign n5468 =  n5452 & ~n5467;
assign n5469 = ~n0019 & ~n0157;
assign n5470 =  n5468 & ~n5469;
assign n5471 =  n0013 & ~n0157;
assign n5472 =  n5470 & ~n5471;
assign n5473 = ~n0022 & ~n0156;
assign n5474 =  n5472 & ~n5473;
assign n5475 = ~n0013 & ~n0156;
assign n5476 =  n5474 & ~n5475;
assign n5477 = ~n0060 & ~n0155;
assign n5478 =  n5476 & ~n5477;
assign n5479 = ~n0014 & ~n0155;
assign n5480 =  n5478 & ~n5479;
assign n5481 = ~n0056 & ~n0154;
assign n5482 =  n5480 & ~n5481;
assign n5483 =  n0014 & ~n0154;
assign n5484 =  n5482 & ~n5483;
assign n5485 = ~n0067 &  n2275;
assign n5486 = ~n0066 &  n5485;
assign n5487 = ~n0065 &  n5486;
assign n5488 = ~n0078 &  n5487;
assign n5489 = ~n0072 &  n5488;
assign n5490 = ~n0042 &  n5489;
assign n5491 =  n0098 &  n5490;
assign n5492 =  n0151 &  n5491;
assign n5493 =  n0150 &  n5492;
assign n5494 =  n0096 &  n5493;
assign n5495 =  n0149 &  n5494;
assign n5496 =  n0093 &  n5495;
assign n5497 =  n0092 &  n5496;
assign n5498 = ~n0153 &  n5497;
assign n5499 =  n5484 & ~n5498;
assign n5500 = ~n0020 & ~n0152;
assign n5501 =  n5499 & ~n5500;
assign n5502 = ~n0013 & ~n0152;
assign n5503 =  n5501 & ~n5502;
assign n5504 = ~n0018 & ~n0151;
assign n5505 =  n5503 & ~n5504;
assign n5506 =  n0013 & ~n0151;
assign n5507 =  n5505 & ~n5506;
assign n5508 = ~n0043 & ~n0150;
assign n5509 =  n5507 & ~n5508;
assign n5510 =  n0014 & ~n0150;
assign n5511 =  n5509 & ~n5510;
assign n5512 = ~n0047 & ~n0149;
assign n5513 =  n5511 & ~n5512;
assign n5514 = ~n0014 & ~n0149;
assign n5515 =  n5513 & ~n5514;
assign n5516 = ~n0026 & ~n0029;
assign n5517 =  n0090 &  n5516;
assign n5518 = ~n0064 &  n5517;
assign n5519 = ~n0063 &  n5518;
assign n5520 = ~n0062 &  n5519;
assign n5521 = ~n0077 &  n5520;
assign n5522 = ~n0071 &  n5521;
assign n5523 =  n0147 &  n5522;
assign n5524 =  n0146 &  n5523;
assign n5525 =  n0145 &  n5524;
assign n5526 =  n0087 &  n5525;
assign n5527 =  n0086 &  n5526;
assign n5528 =  n0144 &  n5527;
assign n5529 =  n0083 &  n5528;
assign n5530 = ~n0148 &  n5529;
assign n5531 =  n5515 & ~n5530;
assign n5532 = ~n0034 & ~n0147;
assign n5533 =  n5531 & ~n5532;
assign n5534 = ~n0014 & ~n0147;
assign n5535 =  n5533 & ~n5534;
assign n5536 = ~n0021 & ~n0146;
assign n5537 =  n5535 & ~n5536;
assign n5538 = ~n0013 & ~n0146;
assign n5539 =  n5537 & ~n5538;
assign n5540 = ~n0030 & ~n0145;
assign n5541 =  n5539 & ~n5540;
assign n5542 =  n0014 & ~n0145;
assign n5543 =  n5541 & ~n5542;
assign n5544 = ~n0017 & ~n0144;
assign n5545 =  n5543 & ~n5544;
assign n5546 =  n0013 & ~n0144;
assign n5547 =  n5545 & ~n5546;
assign n5548 =  n0124 & ~n0143;
assign n5549 =  n5547 & ~n5548;
assign n5550 =  n0133 & ~n0143;
assign n5551 =  n5549 & ~n5550;
assign n5552 =  n0142 & ~n0143;
assign n5553 =  n5551 & ~n5552;
assign n5554 = ~n0069 &  n0925;
assign n5555 = ~n0068 &  n5554;
assign n5556 =  n0141 &  n5555;
assign n5557 =  n0140 &  n5556;
assign n5558 =  n0139 &  n5557;
assign n5559 =  n0138 &  n5558;
assign n5560 =  n0137 &  n5559;
assign n5561 =  n0136 &  n5560;
assign n5562 =  n0135 &  n5561;
assign n5563 =  n0134 &  n5562;
assign n5564 = ~n0142 &  n5563;
assign n5565 =  n5553 & ~n5564;
assign n5566 = ~n0061 & ~n0141;
assign n5567 =  n5565 & ~n5566;
assign n5568 = ~n0014 & ~n0141;
assign n5569 =  n5567 & ~n5568;
assign n5570 = ~n0060 & ~n0140;
assign n5571 =  n5569 & ~n5570;
assign n5572 = ~n0010 & ~n0140;
assign n5573 =  n5571 & ~n5572;
assign n5574 = ~n0057 & ~n0139;
assign n5575 =  n5573 & ~n5574;
assign n5576 =  n0013 & ~n0139;
assign n5577 =  n5575 & ~n5576;
assign n5578 = ~n0022 & ~n0138;
assign n5579 =  n5577 & ~n5578;
assign n5580 = ~n0009 & ~n0138;
assign n5581 =  n5579 & ~n5580;
assign n5582 = ~n0019 & ~n0137;
assign n5583 =  n5581 & ~n5582;
assign n5584 =  n0009 & ~n0137;
assign n5585 =  n5583 & ~n5584;
assign n5586 = ~n0059 & ~n0136;
assign n5587 =  n5585 & ~n5586;
assign n5588 = ~n0013 & ~n0136;
assign n5589 =  n5587 & ~n5588;
assign n5590 = ~n0058 & ~n0135;
assign n5591 =  n5589 & ~n5590;
assign n5592 =  n0014 & ~n0135;
assign n5593 =  n5591 & ~n5592;
assign n5594 = ~n0056 & ~n0134;
assign n5595 =  n5593 & ~n5594;
assign n5596 =  n0010 & ~n0134;
assign n5597 =  n5595 & ~n5596;
assign n5598 = ~n0040 &  n5212;
assign n5599 = ~n0065 &  n5598;
assign n5600 = ~n0042 &  n5599;
assign n5601 = ~n0041 &  n5600;
assign n5602 =  n0132 &  n5601;
assign n5603 =  n0131 &  n5602;
assign n5604 =  n0130 &  n5603;
assign n5605 =  n0129 &  n5604;
assign n5606 =  n0128 &  n5605;
assign n5607 =  n0127 &  n5606;
assign n5608 =  n0126 &  n5607;
assign n5609 =  n0125 &  n5608;
assign n5610 = ~n0133 &  n5609;
assign n5611 =  n5597 & ~n5610;
assign n5612 = ~n0020 & ~n0132;
assign n5613 =  n5611 & ~n5612;
assign n5614 = ~n0009 & ~n0132;
assign n5615 =  n5613 & ~n5614;
assign n5616 = ~n0047 & ~n0131;
assign n5617 =  n5615 & ~n5616;
assign n5618 = ~n0010 & ~n0131;
assign n5619 =  n5617 & ~n5618;
assign n5620 = ~n0044 & ~n0130;
assign n5621 =  n5619 & ~n5620;
assign n5622 =  n0013 & ~n0130;
assign n5623 =  n5621 & ~n5622;
assign n5624 = ~n0018 & ~n0129;
assign n5625 =  n5623 & ~n5624;
assign n5626 =  n0009 & ~n0129;
assign n5627 =  n5625 & ~n5626;
assign n5628 = ~n0046 & ~n0128;
assign n5629 =  n5627 & ~n5628;
assign n5630 = ~n0013 & ~n0128;
assign n5631 =  n5629 & ~n5630;
assign n5632 = ~n0043 & ~n0127;
assign n5633 =  n5631 & ~n5632;
assign n5634 =  n0010 & ~n0127;
assign n5635 =  n5633 & ~n5634;
assign n5636 = ~n0048 & ~n0126;
assign n5637 =  n5635 & ~n5636;
assign n5638 = ~n0014 & ~n0126;
assign n5639 =  n5637 & ~n5638;
assign n5640 = ~n0045 & ~n0125;
assign n5641 =  n5639 & ~n5640;
assign n5642 =  n0014 & ~n0125;
assign n5643 =  n5641 & ~n5642;
assign n5644 = ~n0027 &  n5228;
assign n5645 = ~n0026 &  n5644;
assign n5646 = ~n0063 &  n5645;
assign n5647 = ~n0062 &  n5646;
assign n5648 =  n0123 &  n5647;
assign n5649 =  n0122 &  n5648;
assign n5650 =  n0121 &  n5649;
assign n5651 =  n0120 &  n5650;
assign n5652 =  n0119 &  n5651;
assign n5653 =  n0118 &  n5652;
assign n5654 =  n0117 &  n5653;
assign n5655 =  n0116 &  n5654;
assign n5656 = ~n0124 &  n5655;
assign n5657 =  n5643 & ~n5656;
assign n5658 = ~n0021 & ~n0123;
assign n5659 =  n5657 & ~n5658;
assign n5660 = ~n0009 & ~n0123;
assign n5661 =  n5659 & ~n5660;
assign n5662 = ~n0031 & ~n0122;
assign n5663 =  n5661 & ~n5662;
assign n5664 =  n0013 & ~n0122;
assign n5665 =  n5663 & ~n5664;
assign n5666 = ~n0034 & ~n0121;
assign n5667 =  n5665 & ~n5666;
assign n5668 = ~n0010 & ~n0121;
assign n5669 =  n5667 & ~n5668;
assign n5670 = ~n0017 & ~n0120;
assign n5671 =  n5669 & ~n5670;
assign n5672 =  n0009 & ~n0120;
assign n5673 =  n5671 & ~n5672;
assign n5674 = ~n0035 & ~n0119;
assign n5675 =  n5673 & ~n5674;
assign n5676 = ~n0014 & ~n0119;
assign n5677 =  n5675 & ~n5676;
assign n5678 = ~n0033 & ~n0118;
assign n5679 =  n5677 & ~n5678;
assign n5680 = ~n0013 & ~n0118;
assign n5681 =  n5679 & ~n5680;
assign n5682 = ~n0032 & ~n0117;
assign n5683 =  n5681 & ~n5682;
assign n5684 =  n0014 & ~n0117;
assign n5685 =  n5683 & ~n5684;
assign n5686 = ~n0030 & ~n0116;
assign n5687 =  n5685 & ~n5686;
assign n5688 =  n0010 & ~n0116;
assign n5689 =  n5687 & ~n5688;
assign n5690 =  n0110 &  n0912;
assign n5691 = ~n0115 &  n5690;
assign n5692 =  n5689 & ~n5691;
assign n5693 = ~n0018 & ~n0114;
assign n5694 =  n5692 & ~n5693;
assign n5695 =  n0017 & ~n0114;
assign n5696 =  n5694 & ~n5695;
assign n5697 = ~n0021 & ~n0113;
assign n5698 =  n5696 & ~n5697;
assign n5699 =  n0020 & ~n0113;
assign n5700 =  n5698 & ~n5699;
assign n5701 = ~n0019 & ~n0112;
assign n5702 =  n5700 & ~n5701;
assign n5703 =  n0018 & ~n0112;
assign n5704 =  n5702 & ~n5703;
assign n5705 = ~n0020 & ~n0111;
assign n5706 =  n5704 & ~n5705;
assign n5707 =  n0022 & ~n0111;
assign n5708 =  n5706 & ~n5707;
assign n5709 =  n0091 & ~n0110;
assign n5710 =  n5708 & ~n5709;
assign n5711 =  n0100 & ~n0110;
assign n5712 =  n5710 & ~n5711;
assign n5713 =  n0109 & ~n0110;
assign n5714 =  n5712 & ~n5713;
assign n5715 = ~n0069 &  n5195;
assign n5716 = ~n0049 &  n5715;
assign n5717 = ~n0079 &  n5716;
assign n5718 = ~n0073 &  n5717;
assign n5719 = ~n0082 &  n5718;
assign n5720 =  n0108 &  n5719;
assign n5721 =  n0107 &  n5720;
assign n5722 =  n0106 &  n5721;
assign n5723 =  n0105 &  n5722;
assign n5724 =  n0104 &  n5723;
assign n5725 =  n0103 &  n5724;
assign n5726 =  n0102 &  n5725;
assign n5727 =  n0101 &  n5726;
assign n5728 = ~n0109 &  n5727;
assign n5729 =  n5714 & ~n5728;
assign n5730 = ~n0061 & ~n0108;
assign n5731 =  n5729 & ~n5730;
assign n5732 = ~n0016 & ~n0108;
assign n5733 =  n5731 & ~n5732;
assign n5734 = ~n0015 & ~n0107;
assign n5735 =  n5733 & ~n5734;
assign n5736 = ~n0022 & ~n0107;
assign n5737 =  n5735 & ~n5736;
assign n5738 = ~n0060 & ~n0106;
assign n5739 =  n5737 & ~n5738;
assign n5740 = ~n0016 & ~n0106;
assign n5741 =  n5739 & ~n5740;
assign n5742 = ~n0056 & ~n0105;
assign n5743 =  n5741 & ~n5742;
assign n5744 =  n0016 & ~n0105;
assign n5745 =  n5743 & ~n5744;
assign n5746 = ~n0058 & ~n0104;
assign n5747 =  n5745 & ~n5746;
assign n5748 =  n0016 & ~n0104;
assign n5749 =  n5747 & ~n5748;
assign n5750 = ~n0019 & ~n0103;
assign n5751 =  n5749 & ~n5750;
assign n5752 =  n0015 & ~n0103;
assign n5753 =  n5751 & ~n5752;
assign n5754 = ~n0057 & ~n0102;
assign n5755 =  n5753 & ~n5754;
assign n5756 =  n0015 & ~n0102;
assign n5757 =  n5755 & ~n5756;
assign n5758 = ~n0059 & ~n0101;
assign n5759 =  n5757 & ~n5758;
assign n5760 = ~n0015 & ~n0101;
assign n5761 =  n5759 & ~n5760;
assign n5762 = ~n0036 & ~n0081;
assign n5763 = ~n0066 &  n5762;
assign n5764 = ~n0078 &  n5763;
assign n5765 = ~n0072 &  n5764;
assign n5766 = ~n0042 &  n5765;
assign n5767 =  n0099 &  n5766;
assign n5768 = ~n0041 &  n5767;
assign n5769 =  n0098 &  n5768;
assign n5770 =  n0097 &  n5769;
assign n5771 =  n0096 &  n5770;
assign n5772 =  n0095 &  n5771;
assign n5773 =  n0094 &  n5772;
assign n5774 =  n0093 &  n5773;
assign n5775 =  n0092 &  n5774;
assign n5776 = ~n0100 &  n5775;
assign n5777 =  n5761 & ~n5776;
assign n5778 = ~n0043 & ~n0099;
assign n5779 =  n5777 & ~n5778;
assign n5780 =  n0016 & ~n0099;
assign n5781 =  n5779 & ~n5780;
assign n5782 = ~n0048 & ~n0098;
assign n5783 =  n5781 & ~n5782;
assign n5784 = ~n0016 & ~n0098;
assign n5785 =  n5783 & ~n5784;
assign n5786 = ~n0047 & ~n0097;
assign n5787 =  n5785 & ~n5786;
assign n5788 = ~n0016 & ~n0097;
assign n5789 =  n5787 & ~n5788;
assign n5790 = ~n0045 & ~n0096;
assign n5791 =  n5789 & ~n5790;
assign n5792 =  n0016 & ~n0096;
assign n5793 =  n5791 & ~n5792;
assign n5794 = ~n0015 & ~n0095;
assign n5795 =  n5793 & ~n5794;
assign n5796 = ~n0020 & ~n0095;
assign n5797 =  n5795 & ~n5796;
assign n5798 = ~n0018 & ~n0094;
assign n5799 =  n5797 & ~n5798;
assign n5800 =  n0015 & ~n0094;
assign n5801 =  n5799 & ~n5800;
assign n5802 = ~n0044 & ~n0093;
assign n5803 =  n5801 & ~n5802;
assign n5804 =  n0015 & ~n0093;
assign n5805 =  n5803 & ~n5804;
assign n5806 = ~n0046 & ~n0092;
assign n5807 =  n5805 & ~n5806;
assign n5808 = ~n0015 & ~n0092;
assign n5809 =  n5807 & ~n5808;
assign n5810 =  n0090 &  n1573;
assign n5811 = ~n0063 &  n5810;
assign n5812 = ~n0077 &  n5811;
assign n5813 = ~n0071 &  n5812;
assign n5814 = ~n0080 &  n5813;
assign n5815 =  n0089 &  n5814;
assign n5816 =  n0088 &  n5815;
assign n5817 =  n0087 &  n5816;
assign n5818 =  n0086 &  n5817;
assign n5819 =  n0085 &  n5818;
assign n5820 =  n0084 &  n5819;
assign n5821 =  n0083 &  n5820;
assign n5822 = ~n0091 &  n5821;
assign n5823 =  n5809 & ~n5822;
assign n5824 = ~n0033 & ~n0090;
assign n5825 =  n5823 & ~n5824;
assign n5826 = ~n0015 & ~n0090;
assign n5827 =  n5825 & ~n5826;
assign n5828 = ~n0030 & ~n0089;
assign n5829 =  n5827 & ~n5828;
assign n5830 =  n0016 & ~n0089;
assign n5831 =  n5829 & ~n5830;
assign n5832 = ~n0034 & ~n0088;
assign n5833 =  n5831 & ~n5832;
assign n5834 = ~n0016 & ~n0088;
assign n5835 =  n5833 & ~n5834;
assign n5836 = ~n0035 & ~n0087;
assign n5837 =  n5835 & ~n5836;
assign n5838 = ~n0016 & ~n0087;
assign n5839 =  n5837 & ~n5838;
assign n5840 = ~n0032 & ~n0086;
assign n5841 =  n5839 & ~n5840;
assign n5842 =  n0016 & ~n0086;
assign n5843 =  n5841 & ~n5842;
assign n5844 = ~n0015 & ~n0085;
assign n5845 =  n5843 & ~n5844;
assign n5846 = ~n0021 & ~n0085;
assign n5847 =  n5845 & ~n5846;
assign n5848 = ~n0017 & ~n0084;
assign n5849 =  n5847 & ~n5848;
assign n5850 =  n0015 & ~n0084;
assign n5851 =  n5849 & ~n5850;
assign n5852 = ~n0031 & ~n0083;
assign n5853 =  n5851 & ~n5852;
assign n5854 =  n0015 & ~n0083;
assign n5855 =  n5853 & ~n5854;
assign n0739 =  n5855;
endmodule

