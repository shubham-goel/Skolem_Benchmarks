// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module factorization22_simplified ( i2[21], i2[20], i2[19], i2[18], i2[17], i2[16], i2[15], i2[14], i2[13], i2[12], i2[11], i1[21], i1[20], i1[19], i1[18], i1[17], i1[16], i1[15], i1[14], i1[13], i1[12], i1[11], a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], o_1 );
input i2[21];
input i2[20];
input i2[19];
input i2[18];
input i2[17];
input i2[16];
input i2[15];
input i2[14];
input i2[13];
input i2[12];
input i2[11];
input i1[21];
input i1[20];
input i1[19];
input i1[18];
input i1[17];
input i1[16];
input i1[15];
input i1[14];
input i1[13];
input i1[12];
input i1[11];
input a[0];
input a[1];
input a[2];
input a[3];
input a[4];
input a[5];
input a[6];
input a[7];
input a[8];
input a[9];
input a[10];
input a[11];
input a[12];
input a[13];
input a[14];
input a[15];
input a[16];
input a[17];
input a[18];
input a[19];
input a[20];
input a[21];
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
assign n_1 =  i2[11] &  i1[11];
assign n_2 =  i2[11] &  i1[12];
assign n_3 =  i2[11] &  i1[13];
assign n_4 =  i2[11] &  i1[14];
assign n_5 =  i2[11] &  i1[15];
assign n_6 =  i2[11] &  i1[16];
assign n_7 =  i2[11] &  i1[17];
assign n_8 =  i2[11] &  i1[18];
assign n_9 =  i2[11] &  i1[19];
assign n_10 =  i2[12] &  i1[20];
assign n_11 =  i2[11] &  i1[21];
assign n_12 =  n_10 &  n_11;
assign n_13 =  i2[13] &  i1[20];
assign n_14 =  i2[12] &  i1[21];
assign n_15 =  n_13 &  n_14;
assign n_16 =  i2[14] &  i1[20];
assign n_17 =  i2[13] &  i1[21];
assign n_18 =  n_16 &  n_17;
assign n_19 =  i2[15] &  i1[20];
assign n_20 =  i2[14] &  i1[21];
assign n_21 =  n_19 &  n_20;
assign n_22 =  i2[16] &  i1[20];
assign n_23 =  i2[15] &  i1[21];
assign n_24 =  n_22 &  n_23;
assign n_25 =  i2[17] &  i1[20];
assign n_26 =  i2[16] &  i1[21];
assign n_27 =  n_25 &  n_26;
assign n_28 =  i2[18] &  i1[20];
assign n_29 =  i2[17] &  i1[21];
assign n_30 =  n_28 &  n_29;
assign n_31 =  i2[19] &  i1[20];
assign n_32 =  i2[18] &  i1[21];
assign n_33 =  n_31 &  n_32;
assign n_34 =  i2[20] &  i1[21];
assign n_35 =  i2[21] &  i1[20];
assign n_36 =  n_34 &  n_35;
assign n_37 =  i2[20] &  i1[20];
assign n_38 =  i2[19] &  i1[21];
assign n_39 =  n_37 &  n_38;
assign n_40 = ~n_36 & ~n_39;
assign n_41 = ~n_31 & ~n_32;
assign n_42 = ~n_41 & ~n_33;
assign n_43 = ~n_40 &  n_42;
assign n_44 = ~n_33 & ~n_43;
assign n_45 = ~n_28 & ~n_29;
assign n_46 = ~n_45 & ~n_30;
assign n_47 = ~n_44 &  n_46;
assign n_48 = ~n_30 & ~n_47;
assign n_49 = ~n_25 & ~n_26;
assign n_50 = ~n_49 & ~n_27;
assign n_51 = ~n_48 &  n_50;
assign n_52 = ~n_27 & ~n_51;
assign n_53 = ~n_22 & ~n_23;
assign n_54 = ~n_53 & ~n_24;
assign n_55 = ~n_52 &  n_54;
assign n_56 = ~n_24 & ~n_55;
assign n_57 = ~n_19 & ~n_20;
assign n_58 = ~n_57 & ~n_21;
assign n_59 = ~n_56 &  n_58;
assign n_60 = ~n_21 & ~n_59;
assign n_61 = ~n_16 & ~n_17;
assign n_62 = ~n_61 & ~n_18;
assign n_63 = ~n_60 &  n_62;
assign n_64 = ~n_18 & ~n_63;
assign n_65 = ~n_13 & ~n_14;
assign n_66 = ~n_65 & ~n_15;
assign n_67 = ~n_64 &  n_66;
assign n_68 = ~n_15 & ~n_67;
assign n_69 = ~n_10 & ~n_11;
assign n_70 = ~n_69 & ~n_12;
assign n_71 = ~n_68 &  n_70;
assign n_72 = ~n_12 & ~n_71;
assign n_73 =  i2[11] &  i1[20];
assign n_74 = ~n_72 &  n_73;
assign n_75 =  n_9 &  n_74;
assign n_76 =  i2[12] &  i1[19];
assign n_77 =  n_72 & ~n_73;
assign n_78 = ~n_74 & ~n_77;
assign n_79 =  n_76 &  n_78;
assign n_80 =  n_68 & ~n_70;
assign n_81 = ~n_71 & ~n_80;
assign n_82 =  i2[13] &  i1[19];
assign n_83 =  n_81 &  n_82;
assign n_84 =  n_64 & ~n_66;
assign n_85 = ~n_67 & ~n_84;
assign n_86 =  i2[14] &  i1[19];
assign n_87 =  n_85 &  n_86;
assign n_88 =  n_60 & ~n_62;
assign n_89 = ~n_63 & ~n_88;
assign n_90 =  i2[15] &  i1[19];
assign n_91 =  n_89 &  n_90;
assign n_92 =  n_56 & ~n_58;
assign n_93 = ~n_59 & ~n_92;
assign n_94 =  i2[16] &  i1[19];
assign n_95 =  n_93 &  n_94;
assign n_96 =  n_52 & ~n_54;
assign n_97 = ~n_55 & ~n_96;
assign n_98 =  i2[17] &  i1[19];
assign n_99 =  n_97 &  n_98;
assign n_100 =  n_48 & ~n_50;
assign n_101 = ~n_51 & ~n_100;
assign n_102 =  i2[18] &  i1[19];
assign n_103 =  n_101 &  n_102;
assign n_104 =  n_44 & ~n_46;
assign n_105 = ~n_47 & ~n_104;
assign n_106 =  i2[19] &  i1[19];
assign n_107 =  n_105 &  n_106;
assign n_108 =  n_40 & ~n_42;
assign n_109 = ~n_43 & ~n_108;
assign n_110 =  i2[20] &  i1[19];
assign n_111 =  n_109 &  n_110;
assign n_112 =  i2[21] &  i1[19];
assign n_113 =  n_36 &  n_39;
assign n_114 = ~n_40 & ~n_113;
assign n_115 = ~n_37 & ~n_38;
assign n_116 = ~n_114 & ~n_115;
assign n_117 =  n_112 &  n_116;
assign n_118 = ~n_109 & ~n_110;
assign n_119 = ~n_111 & ~n_118;
assign n_120 =  n_117 &  n_119;
assign n_121 = ~n_111 & ~n_120;
assign n_122 = ~n_105 & ~n_106;
assign n_123 = ~n_107 & ~n_122;
assign n_124 = ~n_121 &  n_123;
assign n_125 = ~n_107 & ~n_124;
assign n_126 = ~n_101 & ~n_102;
assign n_127 = ~n_103 & ~n_126;
assign n_128 = ~n_125 &  n_127;
assign n_129 = ~n_103 & ~n_128;
assign n_130 = ~n_97 & ~n_98;
assign n_131 = ~n_99 & ~n_130;
assign n_132 = ~n_129 &  n_131;
assign n_133 = ~n_99 & ~n_132;
assign n_134 = ~n_93 & ~n_94;
assign n_135 = ~n_95 & ~n_134;
assign n_136 = ~n_133 &  n_135;
assign n_137 = ~n_95 & ~n_136;
assign n_138 = ~n_89 & ~n_90;
assign n_139 = ~n_91 & ~n_138;
assign n_140 = ~n_137 &  n_139;
assign n_141 = ~n_91 & ~n_140;
assign n_142 = ~n_85 & ~n_86;
assign n_143 = ~n_87 & ~n_142;
assign n_144 = ~n_141 &  n_143;
assign n_145 = ~n_87 & ~n_144;
assign n_146 = ~n_81 & ~n_82;
assign n_147 = ~n_83 & ~n_146;
assign n_148 = ~n_145 &  n_147;
assign n_149 = ~n_83 & ~n_148;
assign n_150 = ~n_76 & ~n_78;
assign n_151 = ~n_79 & ~n_150;
assign n_152 = ~n_149 &  n_151;
assign n_153 = ~n_79 & ~n_152;
assign n_154 = ~n_9 & ~n_74;
assign n_155 = ~n_75 & ~n_154;
assign n_156 = ~n_153 &  n_155;
assign n_157 = ~n_75 & ~n_156;
assign n_158 =  n_8 & ~n_157;
assign n_159 =  i2[12] &  i1[18];
assign n_160 =  n_153 & ~n_155;
assign n_161 = ~n_156 & ~n_160;
assign n_162 =  n_159 &  n_161;
assign n_163 =  i2[13] &  i1[18];
assign n_164 =  n_149 & ~n_151;
assign n_165 = ~n_152 & ~n_164;
assign n_166 =  n_163 &  n_165;
assign n_167 =  n_145 & ~n_147;
assign n_168 = ~n_148 & ~n_167;
assign n_169 =  i2[14] &  i1[18];
assign n_170 =  n_168 &  n_169;
assign n_171 =  n_141 & ~n_143;
assign n_172 = ~n_144 & ~n_171;
assign n_173 =  i2[15] &  i1[18];
assign n_174 =  n_172 &  n_173;
assign n_175 =  n_137 & ~n_139;
assign n_176 = ~n_140 & ~n_175;
assign n_177 =  i2[16] &  i1[18];
assign n_178 =  n_176 &  n_177;
assign n_179 =  n_133 & ~n_135;
assign n_180 = ~n_136 & ~n_179;
assign n_181 =  i2[17] &  i1[18];
assign n_182 =  n_180 &  n_181;
assign n_183 =  n_129 & ~n_131;
assign n_184 = ~n_132 & ~n_183;
assign n_185 =  i2[18] &  i1[18];
assign n_186 =  n_184 &  n_185;
assign n_187 =  n_125 & ~n_127;
assign n_188 = ~n_128 & ~n_187;
assign n_189 =  i2[19] &  i1[18];
assign n_190 =  n_188 &  n_189;
assign n_191 =  n_121 & ~n_123;
assign n_192 = ~n_124 & ~n_191;
assign n_193 =  i2[20] &  i1[18];
assign n_194 =  n_192 &  n_193;
assign n_195 = ~n_117 & ~n_119;
assign n_196 = ~n_120 & ~n_195;
assign n_197 =  i2[21] &  i1[18];
assign n_198 =  n_196 &  n_197;
assign n_199 = ~n_192 & ~n_193;
assign n_200 = ~n_194 & ~n_199;
assign n_201 =  n_198 &  n_200;
assign n_202 = ~n_194 & ~n_201;
assign n_203 = ~n_188 & ~n_189;
assign n_204 = ~n_190 & ~n_203;
assign n_205 = ~n_202 &  n_204;
assign n_206 = ~n_190 & ~n_205;
assign n_207 = ~n_184 & ~n_185;
assign n_208 = ~n_186 & ~n_207;
assign n_209 = ~n_206 &  n_208;
assign n_210 = ~n_186 & ~n_209;
assign n_211 = ~n_180 & ~n_181;
assign n_212 = ~n_182 & ~n_211;
assign n_213 = ~n_210 &  n_212;
assign n_214 = ~n_182 & ~n_213;
assign n_215 = ~n_176 & ~n_177;
assign n_216 = ~n_178 & ~n_215;
assign n_217 = ~n_214 &  n_216;
assign n_218 = ~n_178 & ~n_217;
assign n_219 = ~n_172 & ~n_173;
assign n_220 = ~n_174 & ~n_219;
assign n_221 = ~n_218 &  n_220;
assign n_222 = ~n_174 & ~n_221;
assign n_223 = ~n_168 & ~n_169;
assign n_224 = ~n_170 & ~n_223;
assign n_225 = ~n_222 &  n_224;
assign n_226 = ~n_170 & ~n_225;
assign n_227 = ~n_163 & ~n_165;
assign n_228 = ~n_166 & ~n_227;
assign n_229 = ~n_226 &  n_228;
assign n_230 = ~n_166 & ~n_229;
assign n_231 = ~n_159 & ~n_161;
assign n_232 = ~n_162 & ~n_231;
assign n_233 = ~n_230 &  n_232;
assign n_234 = ~n_162 & ~n_233;
assign n_235 = ~n_8 &  n_157;
assign n_236 = ~n_158 & ~n_235;
assign n_237 = ~n_234 &  n_236;
assign n_238 = ~n_158 & ~n_237;
assign n_239 =  n_7 & ~n_238;
assign n_240 =  i2[12] &  i1[17];
assign n_241 =  n_234 & ~n_236;
assign n_242 = ~n_237 & ~n_241;
assign n_243 =  n_240 &  n_242;
assign n_244 =  i2[13] &  i1[17];
assign n_245 =  n_230 & ~n_232;
assign n_246 = ~n_233 & ~n_245;
assign n_247 =  n_244 &  n_246;
assign n_248 =  i2[14] &  i1[17];
assign n_249 =  n_226 & ~n_228;
assign n_250 = ~n_229 & ~n_249;
assign n_251 =  n_248 &  n_250;
assign n_252 =  n_222 & ~n_224;
assign n_253 = ~n_225 & ~n_252;
assign n_254 =  i2[15] &  i1[17];
assign n_255 =  n_253 &  n_254;
assign n_256 =  n_218 & ~n_220;
assign n_257 = ~n_221 & ~n_256;
assign n_258 =  i2[16] &  i1[17];
assign n_259 =  n_257 &  n_258;
assign n_260 =  n_214 & ~n_216;
assign n_261 = ~n_217 & ~n_260;
assign n_262 =  i2[17] &  i1[17];
assign n_263 =  n_261 &  n_262;
assign n_264 =  n_210 & ~n_212;
assign n_265 = ~n_213 & ~n_264;
assign n_266 =  i2[18] &  i1[17];
assign n_267 =  n_265 &  n_266;
assign n_268 =  n_206 & ~n_208;
assign n_269 = ~n_209 & ~n_268;
assign n_270 =  i2[19] &  i1[17];
assign n_271 =  n_269 &  n_270;
assign n_272 =  n_202 & ~n_204;
assign n_273 = ~n_205 & ~n_272;
assign n_274 =  i2[20] &  i1[17];
assign n_275 =  n_273 &  n_274;
assign n_276 = ~n_198 & ~n_200;
assign n_277 = ~n_201 & ~n_276;
assign n_278 =  i2[21] &  i1[17];
assign n_279 =  n_277 &  n_278;
assign n_280 = ~n_273 & ~n_274;
assign n_281 = ~n_275 & ~n_280;
assign n_282 =  n_279 &  n_281;
assign n_283 = ~n_275 & ~n_282;
assign n_284 = ~n_269 & ~n_270;
assign n_285 = ~n_271 & ~n_284;
assign n_286 = ~n_283 &  n_285;
assign n_287 = ~n_271 & ~n_286;
assign n_288 = ~n_265 & ~n_266;
assign n_289 = ~n_267 & ~n_288;
assign n_290 = ~n_287 &  n_289;
assign n_291 = ~n_267 & ~n_290;
assign n_292 = ~n_261 & ~n_262;
assign n_293 = ~n_263 & ~n_292;
assign n_294 = ~n_291 &  n_293;
assign n_295 = ~n_263 & ~n_294;
assign n_296 = ~n_257 & ~n_258;
assign n_297 = ~n_259 & ~n_296;
assign n_298 = ~n_295 &  n_297;
assign n_299 = ~n_259 & ~n_298;
assign n_300 = ~n_253 & ~n_254;
assign n_301 = ~n_255 & ~n_300;
assign n_302 = ~n_299 &  n_301;
assign n_303 = ~n_255 & ~n_302;
assign n_304 = ~n_248 & ~n_250;
assign n_305 = ~n_251 & ~n_304;
assign n_306 = ~n_303 &  n_305;
assign n_307 = ~n_251 & ~n_306;
assign n_308 = ~n_244 & ~n_246;
assign n_309 = ~n_247 & ~n_308;
assign n_310 = ~n_307 &  n_309;
assign n_311 = ~n_247 & ~n_310;
assign n_312 = ~n_240 & ~n_242;
assign n_313 = ~n_243 & ~n_312;
assign n_314 = ~n_311 &  n_313;
assign n_315 = ~n_243 & ~n_314;
assign n_316 = ~n_7 &  n_238;
assign n_317 = ~n_239 & ~n_316;
assign n_318 = ~n_315 &  n_317;
assign n_319 = ~n_239 & ~n_318;
assign n_320 =  n_6 & ~n_319;
assign n_321 =  i2[12] &  i1[16];
assign n_322 =  n_315 & ~n_317;
assign n_323 = ~n_318 & ~n_322;
assign n_324 =  n_321 &  n_323;
assign n_325 =  i2[13] &  i1[16];
assign n_326 =  n_311 & ~n_313;
assign n_327 = ~n_314 & ~n_326;
assign n_328 =  n_325 &  n_327;
assign n_329 =  i2[14] &  i1[16];
assign n_330 =  n_307 & ~n_309;
assign n_331 = ~n_310 & ~n_330;
assign n_332 =  n_329 &  n_331;
assign n_333 =  i2[15] &  i1[16];
assign n_334 =  n_303 & ~n_305;
assign n_335 = ~n_306 & ~n_334;
assign n_336 =  n_333 &  n_335;
assign n_337 =  n_299 & ~n_301;
assign n_338 = ~n_302 & ~n_337;
assign n_339 =  i2[16] &  i1[16];
assign n_340 =  n_338 &  n_339;
assign n_341 =  n_295 & ~n_297;
assign n_342 = ~n_298 & ~n_341;
assign n_343 =  i2[17] &  i1[16];
assign n_344 =  n_342 &  n_343;
assign n_345 =  n_291 & ~n_293;
assign n_346 = ~n_294 & ~n_345;
assign n_347 =  i2[18] &  i1[16];
assign n_348 =  n_346 &  n_347;
assign n_349 =  n_287 & ~n_289;
assign n_350 = ~n_290 & ~n_349;
assign n_351 =  i2[19] &  i1[16];
assign n_352 =  n_350 &  n_351;
assign n_353 =  n_283 & ~n_285;
assign n_354 = ~n_286 & ~n_353;
assign n_355 =  i2[20] &  i1[16];
assign n_356 =  n_354 &  n_355;
assign n_357 = ~n_279 & ~n_281;
assign n_358 = ~n_282 & ~n_357;
assign n_359 =  i2[21] &  i1[16];
assign n_360 =  n_358 &  n_359;
assign n_361 = ~n_354 & ~n_355;
assign n_362 = ~n_356 & ~n_361;
assign n_363 =  n_360 &  n_362;
assign n_364 = ~n_356 & ~n_363;
assign n_365 = ~n_350 & ~n_351;
assign n_366 = ~n_352 & ~n_365;
assign n_367 = ~n_364 &  n_366;
assign n_368 = ~n_352 & ~n_367;
assign n_369 = ~n_346 & ~n_347;
assign n_370 = ~n_348 & ~n_369;
assign n_371 = ~n_368 &  n_370;
assign n_372 = ~n_348 & ~n_371;
assign n_373 = ~n_342 & ~n_343;
assign n_374 = ~n_344 & ~n_373;
assign n_375 = ~n_372 &  n_374;
assign n_376 = ~n_344 & ~n_375;
assign n_377 = ~n_338 & ~n_339;
assign n_378 = ~n_340 & ~n_377;
assign n_379 = ~n_376 &  n_378;
assign n_380 = ~n_340 & ~n_379;
assign n_381 = ~n_333 & ~n_335;
assign n_382 = ~n_336 & ~n_381;
assign n_383 = ~n_380 &  n_382;
assign n_384 = ~n_336 & ~n_383;
assign n_385 = ~n_329 & ~n_331;
assign n_386 = ~n_332 & ~n_385;
assign n_387 = ~n_384 &  n_386;
assign n_388 = ~n_332 & ~n_387;
assign n_389 = ~n_325 & ~n_327;
assign n_390 = ~n_328 & ~n_389;
assign n_391 = ~n_388 &  n_390;
assign n_392 = ~n_328 & ~n_391;
assign n_393 = ~n_321 & ~n_323;
assign n_394 = ~n_324 & ~n_393;
assign n_395 = ~n_392 &  n_394;
assign n_396 = ~n_324 & ~n_395;
assign n_397 = ~n_6 &  n_319;
assign n_398 = ~n_320 & ~n_397;
assign n_399 = ~n_396 &  n_398;
assign n_400 = ~n_320 & ~n_399;
assign n_401 =  n_5 & ~n_400;
assign n_402 =  i2[12] &  i1[15];
assign n_403 =  n_396 & ~n_398;
assign n_404 = ~n_399 & ~n_403;
assign n_405 =  n_402 &  n_404;
assign n_406 =  i2[13] &  i1[15];
assign n_407 =  n_392 & ~n_394;
assign n_408 = ~n_395 & ~n_407;
assign n_409 =  n_406 &  n_408;
assign n_410 =  i2[14] &  i1[15];
assign n_411 =  n_388 & ~n_390;
assign n_412 = ~n_391 & ~n_411;
assign n_413 =  n_410 &  n_412;
assign n_414 =  i2[15] &  i1[15];
assign n_415 =  n_384 & ~n_386;
assign n_416 = ~n_387 & ~n_415;
assign n_417 =  n_414 &  n_416;
assign n_418 =  i2[16] &  i1[15];
assign n_419 =  n_380 & ~n_382;
assign n_420 = ~n_383 & ~n_419;
assign n_421 =  n_418 &  n_420;
assign n_422 =  n_376 & ~n_378;
assign n_423 = ~n_379 & ~n_422;
assign n_424 =  i2[17] &  i1[15];
assign n_425 =  n_423 &  n_424;
assign n_426 =  n_372 & ~n_374;
assign n_427 = ~n_375 & ~n_426;
assign n_428 =  i2[18] &  i1[15];
assign n_429 =  n_427 &  n_428;
assign n_430 =  n_368 & ~n_370;
assign n_431 = ~n_371 & ~n_430;
assign n_432 =  i2[19] &  i1[15];
assign n_433 =  n_431 &  n_432;
assign n_434 =  n_364 & ~n_366;
assign n_435 = ~n_367 & ~n_434;
assign n_436 =  i2[20] &  i1[15];
assign n_437 =  n_435 &  n_436;
assign n_438 = ~n_360 & ~n_362;
assign n_439 = ~n_363 & ~n_438;
assign n_440 =  i2[21] &  i1[15];
assign n_441 =  n_439 &  n_440;
assign n_442 = ~n_435 & ~n_436;
assign n_443 = ~n_437 & ~n_442;
assign n_444 =  n_441 &  n_443;
assign n_445 = ~n_437 & ~n_444;
assign n_446 = ~n_431 & ~n_432;
assign n_447 = ~n_433 & ~n_446;
assign n_448 = ~n_445 &  n_447;
assign n_449 = ~n_433 & ~n_448;
assign n_450 = ~n_427 & ~n_428;
assign n_451 = ~n_429 & ~n_450;
assign n_452 = ~n_449 &  n_451;
assign n_453 = ~n_429 & ~n_452;
assign n_454 = ~n_423 & ~n_424;
assign n_455 = ~n_425 & ~n_454;
assign n_456 = ~n_453 &  n_455;
assign n_457 = ~n_425 & ~n_456;
assign n_458 = ~n_418 & ~n_420;
assign n_459 = ~n_421 & ~n_458;
assign n_460 = ~n_457 &  n_459;
assign n_461 = ~n_421 & ~n_460;
assign n_462 = ~n_414 & ~n_416;
assign n_463 = ~n_417 & ~n_462;
assign n_464 = ~n_461 &  n_463;
assign n_465 = ~n_417 & ~n_464;
assign n_466 = ~n_410 & ~n_412;
assign n_467 = ~n_413 & ~n_466;
assign n_468 = ~n_465 &  n_467;
assign n_469 = ~n_413 & ~n_468;
assign n_470 = ~n_406 & ~n_408;
assign n_471 = ~n_409 & ~n_470;
assign n_472 = ~n_469 &  n_471;
assign n_473 = ~n_409 & ~n_472;
assign n_474 = ~n_402 & ~n_404;
assign n_475 = ~n_405 & ~n_474;
assign n_476 = ~n_473 &  n_475;
assign n_477 = ~n_405 & ~n_476;
assign n_478 = ~n_5 &  n_400;
assign n_479 = ~n_401 & ~n_478;
assign n_480 = ~n_477 &  n_479;
assign n_481 = ~n_401 & ~n_480;
assign n_482 =  n_4 & ~n_481;
assign n_483 =  i2[12] &  i1[14];
assign n_484 =  n_477 & ~n_479;
assign n_485 = ~n_480 & ~n_484;
assign n_486 =  n_483 &  n_485;
assign n_487 =  i2[13] &  i1[14];
assign n_488 =  n_473 & ~n_475;
assign n_489 = ~n_476 & ~n_488;
assign n_490 =  n_487 &  n_489;
assign n_491 =  i2[14] &  i1[14];
assign n_492 =  n_469 & ~n_471;
assign n_493 = ~n_472 & ~n_492;
assign n_494 =  n_491 &  n_493;
assign n_495 =  i2[15] &  i1[14];
assign n_496 =  n_465 & ~n_467;
assign n_497 = ~n_468 & ~n_496;
assign n_498 =  n_495 &  n_497;
assign n_499 =  i2[16] &  i1[14];
assign n_500 =  n_461 & ~n_463;
assign n_501 = ~n_464 & ~n_500;
assign n_502 =  n_499 &  n_501;
assign n_503 =  i2[17] &  i1[14];
assign n_504 =  n_457 & ~n_459;
assign n_505 = ~n_460 & ~n_504;
assign n_506 =  n_503 &  n_505;
assign n_507 =  n_453 & ~n_455;
assign n_508 = ~n_456 & ~n_507;
assign n_509 =  i2[18] &  i1[14];
assign n_510 =  n_508 &  n_509;
assign n_511 =  n_449 & ~n_451;
assign n_512 = ~n_452 & ~n_511;
assign n_513 =  i2[19] &  i1[14];
assign n_514 =  n_512 &  n_513;
assign n_515 =  n_445 & ~n_447;
assign n_516 = ~n_448 & ~n_515;
assign n_517 =  i2[20] &  i1[14];
assign n_518 =  n_516 &  n_517;
assign n_519 = ~n_441 & ~n_443;
assign n_520 = ~n_444 & ~n_519;
assign n_521 =  i2[21] &  i1[14];
assign n_522 =  n_520 &  n_521;
assign n_523 = ~n_516 & ~n_517;
assign n_524 = ~n_518 & ~n_523;
assign n_525 =  n_522 &  n_524;
assign n_526 = ~n_518 & ~n_525;
assign n_527 = ~n_512 & ~n_513;
assign n_528 = ~n_514 & ~n_527;
assign n_529 = ~n_526 &  n_528;
assign n_530 = ~n_514 & ~n_529;
assign n_531 = ~n_508 & ~n_509;
assign n_532 = ~n_510 & ~n_531;
assign n_533 = ~n_530 &  n_532;
assign n_534 = ~n_510 & ~n_533;
assign n_535 = ~n_503 & ~n_505;
assign n_536 = ~n_506 & ~n_535;
assign n_537 = ~n_534 &  n_536;
assign n_538 = ~n_506 & ~n_537;
assign n_539 = ~n_499 & ~n_501;
assign n_540 = ~n_502 & ~n_539;
assign n_541 = ~n_538 &  n_540;
assign n_542 = ~n_502 & ~n_541;
assign n_543 = ~n_495 & ~n_497;
assign n_544 = ~n_498 & ~n_543;
assign n_545 = ~n_542 &  n_544;
assign n_546 = ~n_498 & ~n_545;
assign n_547 = ~n_491 & ~n_493;
assign n_548 = ~n_494 & ~n_547;
assign n_549 = ~n_546 &  n_548;
assign n_550 = ~n_494 & ~n_549;
assign n_551 = ~n_487 & ~n_489;
assign n_552 = ~n_490 & ~n_551;
assign n_553 = ~n_550 &  n_552;
assign n_554 = ~n_490 & ~n_553;
assign n_555 = ~n_483 & ~n_485;
assign n_556 = ~n_486 & ~n_555;
assign n_557 = ~n_554 &  n_556;
assign n_558 = ~n_486 & ~n_557;
assign n_559 = ~n_4 &  n_481;
assign n_560 = ~n_482 & ~n_559;
assign n_561 = ~n_558 &  n_560;
assign n_562 = ~n_482 & ~n_561;
assign n_563 =  n_3 & ~n_562;
assign n_564 =  i2[12] &  i1[13];
assign n_565 =  n_558 & ~n_560;
assign n_566 = ~n_561 & ~n_565;
assign n_567 =  n_564 &  n_566;
assign n_568 =  i2[13] &  i1[13];
assign n_569 =  n_554 & ~n_556;
assign n_570 = ~n_557 & ~n_569;
assign n_571 =  n_568 &  n_570;
assign n_572 =  i2[14] &  i1[13];
assign n_573 =  n_550 & ~n_552;
assign n_574 = ~n_553 & ~n_573;
assign n_575 =  n_572 &  n_574;
assign n_576 =  i2[15] &  i1[13];
assign n_577 =  n_546 & ~n_548;
assign n_578 = ~n_549 & ~n_577;
assign n_579 =  n_576 &  n_578;
assign n_580 =  i2[16] &  i1[13];
assign n_581 =  n_542 & ~n_544;
assign n_582 = ~n_545 & ~n_581;
assign n_583 =  n_580 &  n_582;
assign n_584 =  i2[17] &  i1[13];
assign n_585 =  n_538 & ~n_540;
assign n_586 = ~n_541 & ~n_585;
assign n_587 =  n_584 &  n_586;
assign n_588 =  i2[18] &  i1[13];
assign n_589 =  n_534 & ~n_536;
assign n_590 = ~n_537 & ~n_589;
assign n_591 =  n_588 &  n_590;
assign n_592 =  n_530 & ~n_532;
assign n_593 = ~n_533 & ~n_592;
assign n_594 =  i2[19] &  i1[13];
assign n_595 =  n_593 &  n_594;
assign n_596 =  n_526 & ~n_528;
assign n_597 = ~n_529 & ~n_596;
assign n_598 =  i2[20] &  i1[13];
assign n_599 =  n_597 &  n_598;
assign n_600 = ~n_522 & ~n_524;
assign n_601 = ~n_525 & ~n_600;
assign n_602 =  i2[21] &  i1[13];
assign n_603 =  n_601 &  n_602;
assign n_604 = ~n_597 & ~n_598;
assign n_605 = ~n_599 & ~n_604;
assign n_606 =  n_603 &  n_605;
assign n_607 = ~n_599 & ~n_606;
assign n_608 = ~n_593 & ~n_594;
assign n_609 = ~n_595 & ~n_608;
assign n_610 = ~n_607 &  n_609;
assign n_611 = ~n_595 & ~n_610;
assign n_612 = ~n_588 & ~n_590;
assign n_613 = ~n_591 & ~n_612;
assign n_614 = ~n_611 &  n_613;
assign n_615 = ~n_591 & ~n_614;
assign n_616 = ~n_584 & ~n_586;
assign n_617 = ~n_587 & ~n_616;
assign n_618 = ~n_615 &  n_617;
assign n_619 = ~n_587 & ~n_618;
assign n_620 = ~n_580 & ~n_582;
assign n_621 = ~n_583 & ~n_620;
assign n_622 = ~n_619 &  n_621;
assign n_623 = ~n_583 & ~n_622;
assign n_624 = ~n_576 & ~n_578;
assign n_625 = ~n_579 & ~n_624;
assign n_626 = ~n_623 &  n_625;
assign n_627 = ~n_579 & ~n_626;
assign n_628 = ~n_572 & ~n_574;
assign n_629 = ~n_575 & ~n_628;
assign n_630 = ~n_627 &  n_629;
assign n_631 = ~n_575 & ~n_630;
assign n_632 = ~n_568 & ~n_570;
assign n_633 = ~n_571 & ~n_632;
assign n_634 = ~n_631 &  n_633;
assign n_635 = ~n_571 & ~n_634;
assign n_636 = ~n_564 & ~n_566;
assign n_637 = ~n_567 & ~n_636;
assign n_638 = ~n_635 &  n_637;
assign n_639 = ~n_567 & ~n_638;
assign n_640 = ~n_3 &  n_562;
assign n_641 = ~n_563 & ~n_640;
assign n_642 = ~n_639 &  n_641;
assign n_643 = ~n_563 & ~n_642;
assign n_644 =  n_2 & ~n_643;
assign n_645 =  i2[12] &  i1[12];
assign n_646 =  n_639 & ~n_641;
assign n_647 = ~n_642 & ~n_646;
assign n_648 =  n_645 &  n_647;
assign n_649 =  i2[13] &  i1[12];
assign n_650 =  n_635 & ~n_637;
assign n_651 = ~n_638 & ~n_650;
assign n_652 =  n_649 &  n_651;
assign n_653 =  i2[14] &  i1[12];
assign n_654 =  n_631 & ~n_633;
assign n_655 = ~n_634 & ~n_654;
assign n_656 =  n_653 &  n_655;
assign n_657 =  i2[15] &  i1[12];
assign n_658 =  n_627 & ~n_629;
assign n_659 = ~n_630 & ~n_658;
assign n_660 =  n_657 &  n_659;
assign n_661 =  i2[16] &  i1[12];
assign n_662 =  n_623 & ~n_625;
assign n_663 = ~n_626 & ~n_662;
assign n_664 =  n_661 &  n_663;
assign n_665 =  i2[17] &  i1[12];
assign n_666 =  n_619 & ~n_621;
assign n_667 = ~n_622 & ~n_666;
assign n_668 =  n_665 &  n_667;
assign n_669 =  i2[18] &  i1[12];
assign n_670 =  n_615 & ~n_617;
assign n_671 = ~n_618 & ~n_670;
assign n_672 =  n_669 &  n_671;
assign n_673 =  i2[19] &  i1[12];
assign n_674 =  n_611 & ~n_613;
assign n_675 = ~n_614 & ~n_674;
assign n_676 =  n_673 &  n_675;
assign n_677 =  n_607 & ~n_609;
assign n_678 = ~n_610 & ~n_677;
assign n_679 =  i2[20] &  i1[12];
assign n_680 =  n_678 &  n_679;
assign n_681 = ~n_603 & ~n_605;
assign n_682 = ~n_606 & ~n_681;
assign n_683 =  i2[21] &  i1[12];
assign n_684 =  n_682 &  n_683;
assign n_685 = ~n_678 & ~n_679;
assign n_686 = ~n_680 & ~n_685;
assign n_687 =  n_684 &  n_686;
assign n_688 = ~n_680 & ~n_687;
assign n_689 = ~n_673 & ~n_675;
assign n_690 = ~n_676 & ~n_689;
assign n_691 = ~n_688 &  n_690;
assign n_692 = ~n_676 & ~n_691;
assign n_693 = ~n_669 & ~n_671;
assign n_694 = ~n_672 & ~n_693;
assign n_695 = ~n_692 &  n_694;
assign n_696 = ~n_672 & ~n_695;
assign n_697 = ~n_665 & ~n_667;
assign n_698 = ~n_668 & ~n_697;
assign n_699 = ~n_696 &  n_698;
assign n_700 = ~n_668 & ~n_699;
assign n_701 = ~n_661 & ~n_663;
assign n_702 = ~n_664 & ~n_701;
assign n_703 = ~n_700 &  n_702;
assign n_704 = ~n_664 & ~n_703;
assign n_705 = ~n_657 & ~n_659;
assign n_706 = ~n_660 & ~n_705;
assign n_707 = ~n_704 &  n_706;
assign n_708 = ~n_660 & ~n_707;
assign n_709 = ~n_653 & ~n_655;
assign n_710 = ~n_656 & ~n_709;
assign n_711 = ~n_708 &  n_710;
assign n_712 = ~n_656 & ~n_711;
assign n_713 = ~n_649 & ~n_651;
assign n_714 = ~n_652 & ~n_713;
assign n_715 = ~n_712 &  n_714;
assign n_716 = ~n_652 & ~n_715;
assign n_717 = ~n_645 & ~n_647;
assign n_718 = ~n_648 & ~n_717;
assign n_719 = ~n_716 &  n_718;
assign n_720 = ~n_648 & ~n_719;
assign n_721 = ~n_2 &  n_643;
assign n_722 = ~n_644 & ~n_721;
assign n_723 = ~n_720 &  n_722;
assign n_724 = ~n_644 & ~n_723;
assign n_725 =  n_1 & ~n_724;
assign n_726 =  i2[12] &  i1[11];
assign n_727 =  n_720 & ~n_722;
assign n_728 = ~n_723 & ~n_727;
assign n_729 =  n_726 &  n_728;
assign n_730 =  i2[13] &  i1[11];
assign n_731 =  n_716 & ~n_718;
assign n_732 = ~n_719 & ~n_731;
assign n_733 =  n_730 &  n_732;
assign n_734 =  i2[14] &  i1[11];
assign n_735 =  n_712 & ~n_714;
assign n_736 = ~n_715 & ~n_735;
assign n_737 =  n_734 &  n_736;
assign n_738 =  i2[15] &  i1[11];
assign n_739 =  n_708 & ~n_710;
assign n_740 = ~n_711 & ~n_739;
assign n_741 =  n_738 &  n_740;
assign n_742 =  i2[16] &  i1[11];
assign n_743 =  n_704 & ~n_706;
assign n_744 = ~n_707 & ~n_743;
assign n_745 =  n_742 &  n_744;
assign n_746 =  i2[17] &  i1[11];
assign n_747 =  n_700 & ~n_702;
assign n_748 = ~n_703 & ~n_747;
assign n_749 =  n_746 &  n_748;
assign n_750 =  i2[18] &  i1[11];
assign n_751 =  n_696 & ~n_698;
assign n_752 = ~n_699 & ~n_751;
assign n_753 =  n_750 &  n_752;
assign n_754 =  i2[19] &  i1[11];
assign n_755 =  n_692 & ~n_694;
assign n_756 = ~n_695 & ~n_755;
assign n_757 =  n_754 &  n_756;
assign n_758 =  i2[20] &  i1[11];
assign n_759 =  n_688 & ~n_690;
assign n_760 = ~n_691 & ~n_759;
assign n_761 =  n_758 &  n_760;
assign n_762 = ~n_684 & ~n_686;
assign n_763 = ~n_687 & ~n_762;
assign n_764 =  i2[21] &  i1[11];
assign n_765 =  n_763 &  n_764;
assign n_766 = ~n_758 & ~n_760;
assign n_767 = ~n_761 & ~n_766;
assign n_768 =  n_765 &  n_767;
assign n_769 = ~n_761 & ~n_768;
assign n_770 = ~n_754 & ~n_756;
assign n_771 = ~n_757 & ~n_770;
assign n_772 = ~n_769 &  n_771;
assign n_773 = ~n_757 & ~n_772;
assign n_774 = ~n_750 & ~n_752;
assign n_775 = ~n_753 & ~n_774;
assign n_776 = ~n_773 &  n_775;
assign n_777 = ~n_753 & ~n_776;
assign n_778 = ~n_746 & ~n_748;
assign n_779 = ~n_749 & ~n_778;
assign n_780 = ~n_777 &  n_779;
assign n_781 = ~n_749 & ~n_780;
assign n_782 = ~n_742 & ~n_744;
assign n_783 = ~n_745 & ~n_782;
assign n_784 = ~n_781 &  n_783;
assign n_785 = ~n_745 & ~n_784;
assign n_786 = ~n_738 & ~n_740;
assign n_787 = ~n_741 & ~n_786;
assign n_788 = ~n_785 &  n_787;
assign n_789 = ~n_741 & ~n_788;
assign n_790 = ~n_734 & ~n_736;
assign n_791 = ~n_737 & ~n_790;
assign n_792 = ~n_789 &  n_791;
assign n_793 = ~n_737 & ~n_792;
assign n_794 = ~n_730 & ~n_732;
assign n_795 = ~n_733 & ~n_794;
assign n_796 = ~n_793 &  n_795;
assign n_797 = ~n_733 & ~n_796;
assign n_798 = ~n_726 & ~n_728;
assign n_799 = ~n_729 & ~n_798;
assign n_800 = ~n_797 &  n_799;
assign n_801 = ~n_729 & ~n_800;
assign n_802 = ~n_1 &  n_724;
assign n_803 = ~n_725 & ~n_802;
assign n_804 = ~n_801 &  n_803;
assign n_805 = ~n_725 & ~n_804;
assign n_806 =  a[0] &  n_805;
assign n_807 = ~a[0] & ~n_805;
assign n_808 =  n_801 & ~n_803;
assign n_809 = ~n_804 & ~n_808;
assign n_810 = ~a[1] &  n_809;
assign n_811 =  a[1] & ~n_809;
assign n_812 =  n_797 & ~n_799;
assign n_813 = ~n_800 & ~n_812;
assign n_814 = ~a[2] &  n_813;
assign n_815 =  a[2] & ~n_813;
assign n_816 =  n_793 & ~n_795;
assign n_817 = ~n_796 & ~n_816;
assign n_818 = ~a[3] &  n_817;
assign n_819 =  a[3] & ~n_817;
assign n_820 =  n_789 & ~n_791;
assign n_821 = ~n_792 & ~n_820;
assign n_822 = ~a[4] &  n_821;
assign n_823 =  a[4] & ~n_821;
assign n_824 =  n_785 & ~n_787;
assign n_825 = ~n_788 & ~n_824;
assign n_826 = ~a[5] &  n_825;
assign n_827 =  a[5] & ~n_825;
assign n_828 =  n_781 & ~n_783;
assign n_829 = ~n_784 & ~n_828;
assign n_830 = ~a[6] &  n_829;
assign n_831 =  a[6] & ~n_829;
assign n_832 =  n_777 & ~n_779;
assign n_833 = ~n_780 & ~n_832;
assign n_834 = ~a[7] &  n_833;
assign n_835 =  a[7] & ~n_833;
assign n_836 =  n_773 & ~n_775;
assign n_837 = ~n_776 & ~n_836;
assign n_838 = ~a[8] &  n_837;
assign n_839 =  a[8] & ~n_837;
assign n_840 =  n_769 & ~n_771;
assign n_841 = ~n_772 & ~n_840;
assign n_842 = ~a[9] &  n_841;
assign n_843 =  a[9] & ~n_841;
assign n_844 = ~n_765 & ~n_767;
assign n_845 = ~n_768 & ~n_844;
assign n_846 = ~a[10] &  n_845;
assign n_847 =  a[10] & ~n_845;
assign n_848 = ~n_763 & ~n_764;
assign n_849 = ~n_765 & ~n_848;
assign n_850 = ~a[11] &  n_849;
assign n_851 =  a[11] & ~n_849;
assign n_852 = ~n_682 & ~n_683;
assign n_853 = ~n_684 & ~n_852;
assign n_854 = ~a[12] &  n_853;
assign n_855 =  a[12] & ~n_853;
assign n_856 = ~n_601 & ~n_602;
assign n_857 = ~n_603 & ~n_856;
assign n_858 = ~a[13] &  n_857;
assign n_859 =  a[13] & ~n_857;
assign n_860 = ~n_520 & ~n_521;
assign n_861 = ~n_522 & ~n_860;
assign n_862 = ~a[14] &  n_861;
assign n_863 =  a[14] & ~n_861;
assign n_864 = ~n_439 & ~n_440;
assign n_865 = ~n_441 & ~n_864;
assign n_866 = ~a[15] &  n_865;
assign n_867 =  a[15] & ~n_865;
assign n_868 = ~n_358 & ~n_359;
assign n_869 = ~n_360 & ~n_868;
assign n_870 = ~a[16] &  n_869;
assign n_871 =  a[16] & ~n_869;
assign n_872 = ~n_277 & ~n_278;
assign n_873 = ~n_279 & ~n_872;
assign n_874 = ~a[17] &  n_873;
assign n_875 =  a[17] & ~n_873;
assign n_876 = ~n_196 & ~n_197;
assign n_877 = ~n_198 & ~n_876;
assign n_878 = ~a[18] &  n_877;
assign n_879 =  a[18] & ~n_877;
assign n_880 = ~n_112 & ~n_116;
assign n_881 = ~n_117 & ~n_880;
assign n_882 = ~a[19] &  n_881;
assign n_883 =  a[19] & ~n_881;
assign n_884 = ~n_34 & ~n_35;
assign n_885 = ~n_36 & ~n_884;
assign n_886 = ~a[20] &  n_885;
assign n_887 =  i2[21] &  i1[21];
assign n_888 = ~a[21] & ~n_887;
assign n_889 =  a[21] &  n_887;
assign n_890 = ~n_888 & ~n_889;
assign n_891 =  a[20] & ~n_885;
assign n_892 = ~n_890 & ~n_891;
assign n_893 = ~n_886 &  n_892;
assign n_894 =  i1[21] & ~i1[20];
assign n_895 = ~i1[19] & ~i1[18];
assign n_896 = ~i1[17] & ~i1[16];
assign n_897 =  n_895 &  n_896;
assign n_898 =  n_894 &  n_897;
assign n_899 = ~i1[15] & ~i1[14];
assign n_900 = ~i1[13] & ~i1[12];
assign n_901 =  n_899 &  n_900;
assign n_902 = ~i1[11] &  n_901;
assign n_903 =  n_898 &  n_902;
assign n_904 =  i2[21] & ~i2[20];
assign n_905 = ~i2[19] & ~i2[18];
assign n_906 = ~i2[17] & ~i2[16];
assign n_907 =  n_905 &  n_906;
assign n_908 =  n_904 &  n_907;
assign n_909 = ~i2[15] & ~i2[14];
assign n_910 = ~i2[13] & ~i2[12];
assign n_911 =  n_909 &  n_910;
assign n_912 = ~i2[11] &  n_911;
assign n_913 =  n_908 &  n_912;
assign n_914 = ~n_903 & ~n_913;
assign n_915 =  n_893 &  n_914;
assign n_916 = ~n_883 &  n_915;
assign n_917 = ~n_882 &  n_916;
assign n_918 = ~n_879 &  n_917;
assign n_919 = ~n_878 &  n_918;
assign n_920 = ~n_875 &  n_919;
assign n_921 = ~n_874 &  n_920;
assign n_922 = ~n_871 &  n_921;
assign n_923 = ~n_870 &  n_922;
assign n_924 = ~n_867 &  n_923;
assign n_925 = ~n_866 &  n_924;
assign n_926 = ~n_863 &  n_925;
assign n_927 = ~n_862 &  n_926;
assign n_928 = ~n_859 &  n_927;
assign n_929 = ~n_858 &  n_928;
assign n_930 = ~n_855 &  n_929;
assign n_931 = ~n_854 &  n_930;
assign n_932 = ~n_851 &  n_931;
assign n_933 = ~n_850 &  n_932;
assign n_934 = ~n_847 &  n_933;
assign n_935 = ~n_846 &  n_934;
assign n_936 = ~n_843 &  n_935;
assign n_937 = ~n_842 &  n_936;
assign n_938 = ~n_839 &  n_937;
assign n_939 = ~n_838 &  n_938;
assign n_940 = ~n_835 &  n_939;
assign n_941 = ~n_834 &  n_940;
assign n_942 = ~n_831 &  n_941;
assign n_943 = ~n_830 &  n_942;
assign n_944 = ~n_827 &  n_943;
assign n_945 = ~n_826 &  n_944;
assign n_946 = ~n_823 &  n_945;
assign n_947 = ~n_822 &  n_946;
assign n_948 = ~n_819 &  n_947;
assign n_949 = ~n_818 &  n_948;
assign n_950 = ~n_815 &  n_949;
assign n_951 = ~n_814 &  n_950;
assign n_952 = ~n_811 &  n_951;
assign n_953 = ~n_810 &  n_952;
assign n_954 = ~n_807 &  n_953;
assign n_955 = ~n_806 &  n_954;
assign o_1 =  n_955;
endmodule

